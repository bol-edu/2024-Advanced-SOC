
//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ../td_ccore_solutions/ROM_1i4_1o8_0bc064f669c474330176c941c6dd719bb8_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   f1921061@cad30
//  Generated date: Tue May 28 14:28:42 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i4_1o8_0bc064f669c474330176c941c6dd719bb8
// ------------------------------------------------------------------


module ROM_1i4_1o8_0bc064f669c474330176c941c6dd719bb8 (
  I_1, O_1
);
  input [3:0] I_1;
  output [7:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_8_12_2(8'b11110000, 8'b11100001, 8'b11010010, 8'b11000011, 8'b10110100,
      8'b10100101, 8'b10010110, 8'b10000111, 8'b01111000, 8'b01101001, 8'b01011010,
      8'b01001011, I_1);

  function automatic [7:0] MUX_v_8_12_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [7:0] input_10;
    input [7:0] input_11;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0000 : begin
        result = input_0;
      end
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      4'b1001 : begin
        result = input_9;
      end
      4'b1010 : begin
        result = input_10;
      end
      default : begin
        result = input_11;
      end
    endcase
    MUX_v_8_12_2 = result;
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/ROM_1i4_1o8_6f8a8acefa07ca761551b27c9076176eb8_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   f1921061@cad30
//  Generated date: Tue May 28 14:28:46 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ROM_1i4_1o8_6f8a8acefa07ca761551b27c9076176eb8
// ------------------------------------------------------------------


module ROM_1i4_1o8_6f8a8acefa07ca761551b27c9076176eb8 (
  I_1, O_1
);
  input [3:0] I_1;
  output [7:0] O_1;



  // Interconnect Declarations for Component Instantiations 
  assign O_1 = MUX_v_8_8_2x4x5(8'b01111000, 8'b01101001, 8'b01011010, 8'b01001011,
      8'b10010110, 8'b10000111, I_1[2:0]);

  function automatic [7:0] MUX_v_8_8_2x4x5;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2x4x5 = result;
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   f1921061@cad30
//  Generated date: Wed Jun  5 13:11:28 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module Encrypt_Top_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, INIT_P12_C_0_tr0, AD_P6_C_0_tr0, ADLEN_C_2_tr0,
      ENC_P6_C_0_tr0, PLEN_C_3_tr0, FINAL_P12_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [18:0] fsm_output;
  reg [18:0] fsm_output;
  input INIT_P12_C_0_tr0;
  input AD_P6_C_0_tr0;
  input ADLEN_C_2_tr0;
  input ENC_P6_C_0_tr0;
  input PLEN_C_3_tr0;
  input FINAL_P12_C_0_tr0;


  // FSM State Type Declaration for Encrypt_Top_run_run_fsm_1
  parameter
    main_C_0 = 5'd0,
    INIT_P12_C_0 = 5'd1,
    ADLEN_C_0 = 5'd2,
    ADLEN_C_1 = 5'd3,
    AD_P6_C_0 = 5'd4,
    ADLEN_C_2 = 5'd5,
    main_C_1 = 5'd6,
    main_C_2 = 5'd7,
    main_C_3 = 5'd8,
    PLEN_C_0 = 5'd9,
    PLEN_C_1 = 5'd10,
    ENC_P6_C_0 = 5'd11,
    PLEN_C_2 = 5'd12,
    PLEN_C_3 = 5'd13,
    FINAL_P12_C_0 = 5'd14,
    main_C_4 = 5'd15,
    main_C_5 = 5'd16,
    main_C_6 = 5'd17,
    main_C_7 = 5'd18;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : Encrypt_Top_run_run_fsm_1
    case (state_var)
      INIT_P12_C_0 : begin
        fsm_output = 19'b0000000000000000010;
        if ( INIT_P12_C_0_tr0 ) begin
          state_var_NS = ADLEN_C_0;
        end
        else begin
          state_var_NS = INIT_P12_C_0;
        end
      end
      ADLEN_C_0 : begin
        fsm_output = 19'b0000000000000000100;
        state_var_NS = ADLEN_C_1;
      end
      ADLEN_C_1 : begin
        fsm_output = 19'b0000000000000001000;
        state_var_NS = AD_P6_C_0;
      end
      AD_P6_C_0 : begin
        fsm_output = 19'b0000000000000010000;
        if ( AD_P6_C_0_tr0 ) begin
          state_var_NS = ADLEN_C_2;
        end
        else begin
          state_var_NS = AD_P6_C_0;
        end
      end
      ADLEN_C_2 : begin
        fsm_output = 19'b0000000000000100000;
        if ( ADLEN_C_2_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = ADLEN_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 19'b0000000000001000000;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 19'b0000000000010000000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 19'b0000000000100000000;
        state_var_NS = PLEN_C_0;
      end
      PLEN_C_0 : begin
        fsm_output = 19'b0000000001000000000;
        state_var_NS = PLEN_C_1;
      end
      PLEN_C_1 : begin
        fsm_output = 19'b0000000010000000000;
        state_var_NS = ENC_P6_C_0;
      end
      ENC_P6_C_0 : begin
        fsm_output = 19'b0000000100000000000;
        if ( ENC_P6_C_0_tr0 ) begin
          state_var_NS = PLEN_C_2;
        end
        else begin
          state_var_NS = ENC_P6_C_0;
        end
      end
      PLEN_C_2 : begin
        fsm_output = 19'b0000001000000000000;
        state_var_NS = PLEN_C_3;
      end
      PLEN_C_3 : begin
        fsm_output = 19'b0000010000000000000;
        if ( PLEN_C_3_tr0 ) begin
          state_var_NS = FINAL_P12_C_0;
        end
        else begin
          state_var_NS = PLEN_C_0;
        end
      end
      FINAL_P12_C_0 : begin
        fsm_output = 19'b0000100000000000000;
        if ( FINAL_P12_C_0_tr0 ) begin
          state_var_NS = main_C_4;
        end
        else begin
          state_var_NS = FINAL_P12_C_0;
        end
      end
      main_C_4 : begin
        fsm_output = 19'b0001000000000000000;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 19'b0010000000000000000;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 19'b0100000000000000000;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 19'b1000000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 19'b0000000000000000001;
        state_var_NS = INIT_P12_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_staller
// ------------------------------------------------------------------


module Encrypt_Top_run_staller (
  run_wen, data_in_rsci_wen_comp, data_out_rsci_wen_comp
);
  output run_wen;
  input data_in_rsci_wen_comp;
  input data_out_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = data_in_rsci_wen_comp & data_out_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_out_rsci_data_out_wait_dp
// ------------------------------------------------------------------


module Encrypt_Top_run_data_out_rsci_data_out_wait_dp (
  clk, rst, arst_n, data_out_rsci_oswt, data_out_rsci_wen_comp, data_out_rsci_biwt,
      data_out_rsci_bdwt, data_out_rsci_bcwt
);
  input clk;
  input rst;
  input arst_n;
  input data_out_rsci_oswt;
  output data_out_rsci_wen_comp;
  input data_out_rsci_biwt;
  input data_out_rsci_bdwt;
  output data_out_rsci_bcwt;
  reg data_out_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign data_out_rsci_wen_comp = (~ data_out_rsci_oswt) | data_out_rsci_biwt | data_out_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      data_out_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      data_out_rsci_bcwt <= 1'b0;
    end
    else begin
      data_out_rsci_bcwt <= ~((~(data_out_rsci_bcwt | data_out_rsci_biwt)) | data_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_out_rsci_data_out_wait_ctrl
// ------------------------------------------------------------------


module Encrypt_Top_run_data_out_rsci_data_out_wait_ctrl (
  run_wen, data_out_rsci_oswt, data_out_rsci_biwt, data_out_rsci_bdwt, data_out_rsci_bcwt,
      data_out_rsci_irdy, data_out_rsci_ivld_run_sct
);
  input run_wen;
  input data_out_rsci_oswt;
  output data_out_rsci_biwt;
  output data_out_rsci_bdwt;
  input data_out_rsci_bcwt;
  input data_out_rsci_irdy;
  output data_out_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire data_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign data_out_rsci_bdwt = data_out_rsci_oswt & run_wen;
  assign data_out_rsci_biwt = data_out_rsci_ogwt & data_out_rsci_irdy;
  assign data_out_rsci_ogwt = data_out_rsci_oswt & (~ data_out_rsci_bcwt);
  assign data_out_rsci_ivld_run_sct = data_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_in_rsci_data_in_wait_dp
// ------------------------------------------------------------------


module Encrypt_Top_run_data_in_rsci_data_in_wait_dp (
  clk, rst, arst_n, data_in_rsci_oswt, data_in_rsci_wen_comp, data_in_rsci_idat_mxwt,
      data_in_rsci_biwt, data_in_rsci_bdwt, data_in_rsci_bcwt, data_in_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  input data_in_rsci_oswt;
  output data_in_rsci_wen_comp;
  output [31:0] data_in_rsci_idat_mxwt;
  input data_in_rsci_biwt;
  input data_in_rsci_bdwt;
  output data_in_rsci_bcwt;
  reg data_in_rsci_bcwt;
  input [31:0] data_in_rsci_idat;


  // Interconnect Declarations
  reg [31:0] data_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign data_in_rsci_wen_comp = (~ data_in_rsci_oswt) | data_in_rsci_biwt | data_in_rsci_bcwt;
  assign data_in_rsci_idat_mxwt = MUX_v_32_2_2(data_in_rsci_idat, data_in_rsci_idat_bfwt,
      data_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      data_in_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      data_in_rsci_bcwt <= 1'b0;
    end
    else begin
      data_in_rsci_bcwt <= ~((~(data_in_rsci_bcwt | data_in_rsci_biwt)) | data_in_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      data_in_rsci_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      data_in_rsci_idat_bfwt <= 32'b00000000000000000000000000000000;
    end
    else if ( data_in_rsci_biwt ) begin
      data_in_rsci_idat_bfwt <= data_in_rsci_idat;
    end
  end

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_in_rsci_data_in_wait_ctrl
// ------------------------------------------------------------------


module Encrypt_Top_run_data_in_rsci_data_in_wait_ctrl (
  run_wen, data_in_rsci_oswt, data_in_rsci_biwt, data_in_rsci_bdwt, data_in_rsci_bcwt,
      data_in_rsci_irdy_run_sct, data_in_rsci_ivld
);
  input run_wen;
  input data_in_rsci_oswt;
  output data_in_rsci_biwt;
  output data_in_rsci_bdwt;
  input data_in_rsci_bcwt;
  output data_in_rsci_irdy_run_sct;
  input data_in_rsci_ivld;


  // Interconnect Declarations
  wire data_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign data_in_rsci_bdwt = data_in_rsci_oswt & run_wen;
  assign data_in_rsci_biwt = data_in_rsci_ogwt & data_in_rsci_ivld;
  assign data_in_rsci_ogwt = data_in_rsci_oswt & (~ data_in_rsci_bcwt);
  assign data_in_rsci_irdy_run_sct = data_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_out_rsci
// ------------------------------------------------------------------


module Encrypt_Top_run_data_out_rsci (
  clk, rst, arst_n, data_out_rsc_dat, data_out_rsc_vld, data_out_rsc_rdy, run_wen,
      data_out_rsci_oswt, data_out_rsci_wen_comp, data_out_rsci_idat
);
  input clk;
  input rst;
  input arst_n;
  output [31:0] data_out_rsc_dat;
  output data_out_rsc_vld;
  input data_out_rsc_rdy;
  input run_wen;
  input data_out_rsci_oswt;
  output data_out_rsci_wen_comp;
  input [31:0] data_out_rsci_idat;


  // Interconnect Declarations
  wire data_out_rsci_biwt;
  wire data_out_rsci_bdwt;
  wire data_out_rsci_bcwt;
  wire data_out_rsci_irdy;
  wire data_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd12),
  .width(32'sd32)) data_out_rsci (
      .irdy(data_out_rsci_irdy),
      .ivld(data_out_rsci_ivld_run_sct),
      .idat(data_out_rsci_idat),
      .rdy(data_out_rsc_rdy),
      .vld(data_out_rsc_vld),
      .dat(data_out_rsc_dat)
    );
  Encrypt_Top_run_data_out_rsci_data_out_wait_ctrl Encrypt_Top_run_data_out_rsci_data_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .data_out_rsci_oswt(data_out_rsci_oswt),
      .data_out_rsci_biwt(data_out_rsci_biwt),
      .data_out_rsci_bdwt(data_out_rsci_bdwt),
      .data_out_rsci_bcwt(data_out_rsci_bcwt),
      .data_out_rsci_irdy(data_out_rsci_irdy),
      .data_out_rsci_ivld_run_sct(data_out_rsci_ivld_run_sct)
    );
  Encrypt_Top_run_data_out_rsci_data_out_wait_dp Encrypt_Top_run_data_out_rsci_data_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .data_out_rsci_oswt(data_out_rsci_oswt),
      .data_out_rsci_wen_comp(data_out_rsci_wen_comp),
      .data_out_rsci_biwt(data_out_rsci_biwt),
      .data_out_rsci_bdwt(data_out_rsci_bdwt),
      .data_out_rsci_bcwt(data_out_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run_data_in_rsci
// ------------------------------------------------------------------


module Encrypt_Top_run_data_in_rsci (
  clk, rst, arst_n, data_in_rsc_dat, data_in_rsc_vld, data_in_rsc_rdy, run_wen, data_in_rsci_oswt,
      data_in_rsci_wen_comp, data_in_rsci_idat_mxwt
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] data_in_rsc_dat;
  input data_in_rsc_vld;
  output data_in_rsc_rdy;
  input run_wen;
  input data_in_rsci_oswt;
  output data_in_rsci_wen_comp;
  output [31:0] data_in_rsci_idat_mxwt;


  // Interconnect Declarations
  wire data_in_rsci_biwt;
  wire data_in_rsci_bdwt;
  wire data_in_rsci_bcwt;
  wire data_in_rsci_irdy_run_sct;
  wire data_in_rsci_ivld;
  wire [31:0] data_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd11),
  .width(32'sd32)) data_in_rsci (
      .rdy(data_in_rsc_rdy),
      .vld(data_in_rsc_vld),
      .dat(data_in_rsc_dat),
      .irdy(data_in_rsci_irdy_run_sct),
      .ivld(data_in_rsci_ivld),
      .idat(data_in_rsci_idat)
    );
  Encrypt_Top_run_data_in_rsci_data_in_wait_ctrl Encrypt_Top_run_data_in_rsci_data_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .data_in_rsci_oswt(data_in_rsci_oswt),
      .data_in_rsci_biwt(data_in_rsci_biwt),
      .data_in_rsci_bdwt(data_in_rsci_bdwt),
      .data_in_rsci_bcwt(data_in_rsci_bcwt),
      .data_in_rsci_irdy_run_sct(data_in_rsci_irdy_run_sct),
      .data_in_rsci_ivld(data_in_rsci_ivld)
    );
  Encrypt_Top_run_data_in_rsci_data_in_wait_dp Encrypt_Top_run_data_in_rsci_data_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .data_in_rsci_oswt(data_in_rsci_oswt),
      .data_in_rsci_wen_comp(data_in_rsci_wen_comp),
      .data_in_rsci_idat_mxwt(data_in_rsci_idat_mxwt),
      .data_in_rsci_biwt(data_in_rsci_biwt),
      .data_in_rsci_bdwt(data_in_rsci_bdwt),
      .data_in_rsci_bcwt(data_in_rsci_bcwt),
      .data_in_rsci_idat(data_in_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top_run
// ------------------------------------------------------------------


module Encrypt_Top_run (
  clk, rst, arst_n, key1, key2, key3, key4, nonce1, nonce2, nonce3, nonce4, adlen,
      plen, data_in_rsc_dat, data_in_rsc_vld, data_in_rsc_rdy, data_out_rsc_dat,
      data_out_rsc_vld, data_out_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] key1;
  input [31:0] key2;
  input [31:0] key3;
  input [31:0] key4;
  input [31:0] nonce1;
  input [31:0] nonce2;
  input [31:0] nonce3;
  input [31:0] nonce4;
  input [7:0] adlen;
  input [7:0] plen;
  input [31:0] data_in_rsc_dat;
  input data_in_rsc_vld;
  output data_in_rsc_rdy;
  output [31:0] data_out_rsc_dat;
  output data_out_rsc_vld;
  input data_out_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire data_in_rsci_wen_comp;
  wire [31:0] data_in_rsci_idat_mxwt;
  wire data_out_rsci_wen_comp;
  reg data_out_rsci_idat_31;
  reg data_out_rsci_idat_30;
  reg data_out_rsci_idat_29;
  reg data_out_rsci_idat_28;
  reg data_out_rsci_idat_27;
  reg data_out_rsci_idat_26;
  reg data_out_rsci_idat_25;
  reg data_out_rsci_idat_24;
  reg data_out_rsci_idat_23;
  reg data_out_rsci_idat_22;
  reg data_out_rsci_idat_21;
  reg data_out_rsci_idat_20;
  reg data_out_rsci_idat_19;
  reg data_out_rsci_idat_18;
  reg data_out_rsci_idat_17;
  reg data_out_rsci_idat_16;
  reg data_out_rsci_idat_15;
  reg data_out_rsci_idat_14;
  reg data_out_rsci_idat_13;
  reg data_out_rsci_idat_12;
  reg data_out_rsci_idat_11;
  reg data_out_rsci_idat_10;
  reg data_out_rsci_idat_9;
  reg data_out_rsci_idat_8;
  reg data_out_rsci_idat_7;
  reg data_out_rsci_idat_6;
  reg data_out_rsci_idat_5;
  reg data_out_rsci_idat_4;
  reg data_out_rsci_idat_3;
  reg data_out_rsci_idat_2;
  reg data_out_rsci_idat_1;
  reg data_out_rsci_idat_0;
  wire [18:0] fsm_output;
  wire operator_33_true_1_operator_33_true_1_and_tmp;
  wire or_dcpl_9;
  wire or_tmp_382;
  wire or_tmp_913;
  wire or_tmp_1693;
  wire and_24_cse;
  wire and_90_cse;
  wire and_94_cse;
  wire and_738_cse;
  wire and_740_cse;
  wire and_885_cse;
  wire and_4636_cse;
  wire xor_2168_cse;
  wire xor_2162_cse;
  wire xor_2172_cse;
  wire xor_2186_cse;
  wire xor_2182_cse;
  wire xor_2184_cse;
  reg reg_data_out_rsci_iswt0_cse;
  reg reg_data_in_rsci_iswt0_cse;
  wire state_and_cse;
  wire state_and_4_cse;
  wire state_and_8_cse;
  wire state_and_24_cse;
  wire state_and_56_cse;
  wire state_and_64_cse;
  wire state_and_86_cse;
  wire state_and_90_cse;
  wire state_and_92_cse;
  wire state_and_98_cse;
  wire state_and_118_cse;
  wire state_and_120_cse;
  wire state_and_128_cse;
  wire state_and_137_cse;
  wire state_and_158_cse;
  wire state_and_161_cse;
  wire state_and_192_cse;
  wire state_and_201_cse;
  wire state_and_208_cse;
  wire and_21_cse;
  wire and_39_cse;
  wire ADLEN_i_and_ssc;
  wire [8:0] z_out;
  wire [9:0] nl_z_out;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  reg state_2_0_1_lpi_4;
  reg state_2_1_1_lpi_4;
  reg state_2_2_1_lpi_4;
  reg state_2_3_1_lpi_4;
  reg state_2_4_1_lpi_4;
  reg state_2_5_1_lpi_4;
  reg state_2_6_1_lpi_4;
  reg state_2_7_1_lpi_4;
  reg state_2_8_1_lpi_4;
  reg state_2_9_1_lpi_4;
  reg state_2_10_1_lpi_4;
  reg state_2_11_1_lpi_4;
  reg state_2_12_1_lpi_4;
  reg state_2_13_1_lpi_4;
  reg state_2_14_1_lpi_4;
  reg state_2_15_1_lpi_4;
  reg state_2_16_1_lpi_4;
  reg state_2_17_1_lpi_4;
  reg state_2_18_1_lpi_4;
  reg state_2_19_1_lpi_4;
  reg state_2_20_1_lpi_4;
  reg state_2_21_1_lpi_4;
  reg state_2_22_1_lpi_4;
  reg state_2_23_1_lpi_4;
  reg state_2_24_1_lpi_4;
  reg state_2_25_1_lpi_4;
  reg state_2_26_1_lpi_4;
  reg state_2_27_1_lpi_4;
  reg state_2_28_1_lpi_4;
  reg state_2_29_1_lpi_4;
  reg state_2_30_1_lpi_4;
  reg state_2_31_1_lpi_4;
  reg state_2_32_1_lpi_4;
  reg state_2_33_1_lpi_4;
  reg state_2_34_1_lpi_4;
  reg state_2_35_1_lpi_4;
  reg state_2_36_1_lpi_4;
  reg state_2_37_1_lpi_4;
  reg state_2_38_1_lpi_4;
  reg state_2_39_1_lpi_4;
  reg state_2_40_1_lpi_4;
  reg state_2_41_1_lpi_4;
  reg state_2_42_1_lpi_4;
  reg state_2_43_1_lpi_4;
  reg state_2_44_1_lpi_4;
  reg state_2_45_1_lpi_4;
  reg state_2_46_1_lpi_4;
  reg state_2_47_1_lpi_4;
  reg state_2_48_1_lpi_4;
  reg state_2_49_1_lpi_4;
  reg state_2_50_1_lpi_4;
  reg state_2_51_1_lpi_4;
  reg state_2_52_1_lpi_4;
  reg state_2_53_1_lpi_4;
  reg state_2_54_1_lpi_4;
  reg state_2_55_1_lpi_4;
  reg state_2_56_1_lpi_4;
  reg state_2_57_1_lpi_4;
  reg state_2_58_1_lpi_4;
  reg state_2_59_1_lpi_4;
  reg state_2_60_1_lpi_4;
  reg state_2_61_1_lpi_4;
  reg state_2_62_1_lpi_4;
  reg state_2_63_1_lpi_4;
  reg state_3_31_lpi_3;
  reg state_3_32_lpi_3;
  reg state_3_30_lpi_3;
  reg state_3_33_lpi_3;
  reg state_3_29_lpi_3;
  reg state_3_34_lpi_3;
  reg state_3_28_lpi_3;
  reg state_3_35_lpi_3;
  reg state_3_27_lpi_3;
  reg state_3_36_lpi_3;
  reg state_3_26_lpi_3;
  reg state_3_37_lpi_3;
  reg state_3_25_lpi_3;
  reg state_3_38_lpi_3;
  reg state_3_24_lpi_3;
  reg state_3_39_lpi_3;
  reg state_3_23_lpi_3;
  reg state_3_40_lpi_3;
  reg state_3_22_lpi_3;
  reg state_3_41_lpi_3;
  reg state_3_21_lpi_3;
  reg state_3_42_lpi_3;
  reg state_3_20_lpi_3;
  reg state_3_43_lpi_3;
  reg state_3_19_lpi_3;
  reg state_3_44_lpi_3;
  reg state_3_18_lpi_3;
  reg state_3_45_lpi_3;
  reg state_3_17_lpi_3;
  reg state_3_46_lpi_3;
  reg state_3_16_lpi_3;
  reg state_3_47_lpi_3;
  reg state_3_15_lpi_3;
  reg state_3_48_lpi_3;
  reg state_3_14_lpi_3;
  reg state_3_49_lpi_3;
  reg state_3_13_lpi_3;
  reg state_3_50_lpi_3;
  reg state_3_12_lpi_3;
  reg state_3_51_lpi_3;
  reg state_3_11_lpi_3;
  reg state_3_52_lpi_3;
  reg state_3_10_lpi_3;
  reg state_3_53_lpi_3;
  reg state_3_9_lpi_3;
  reg state_3_54_lpi_3;
  reg state_3_8_lpi_3;
  reg state_3_55_lpi_3;
  reg state_3_7_lpi_3;
  reg state_3_56_lpi_3;
  reg state_3_6_lpi_3;
  reg state_3_57_lpi_3;
  reg state_3_5_lpi_3;
  reg state_3_58_lpi_3;
  reg state_3_4_lpi_3;
  reg state_3_59_lpi_3;
  reg state_3_3_lpi_3;
  reg state_3_60_lpi_3;
  reg state_3_2_lpi_3;
  reg state_3_61_lpi_3;
  reg state_3_1_lpi_3;
  reg state_3_62_lpi_3;
  reg state_3_0_lpi_3;
  reg state_3_63_lpi_3;
  reg state_4_4_31_lpi_3;
  reg state_4_4_32_lpi_3;
  reg state_4_4_30_lpi_3;
  reg state_4_4_33_lpi_3;
  reg state_4_4_29_lpi_3;
  reg state_4_4_34_lpi_3;
  reg state_4_4_28_lpi_3;
  reg state_4_4_35_lpi_3;
  reg state_4_4_27_lpi_3;
  reg state_4_4_36_lpi_3;
  reg state_4_4_26_lpi_3;
  reg state_4_4_37_lpi_3;
  reg state_4_4_25_lpi_3;
  reg state_4_4_38_lpi_3;
  reg state_4_4_24_lpi_3;
  reg state_4_4_39_lpi_3;
  reg state_4_4_23_lpi_3;
  reg state_4_4_40_lpi_3;
  reg state_4_4_22_lpi_3;
  reg state_4_4_41_lpi_3;
  reg state_4_4_21_lpi_3;
  reg state_4_4_42_lpi_3;
  reg state_4_4_20_lpi_3;
  reg state_4_4_43_lpi_3;
  reg state_4_4_19_lpi_3;
  reg state_4_4_44_lpi_3;
  reg state_4_4_18_lpi_3;
  reg state_4_4_45_lpi_3;
  reg state_4_4_17_lpi_3;
  reg state_4_4_46_lpi_3;
  reg state_4_4_16_lpi_3;
  reg state_4_4_47_lpi_3;
  reg state_4_4_15_lpi_3;
  reg state_4_4_48_lpi_3;
  reg state_4_4_14_lpi_3;
  reg state_4_4_49_lpi_3;
  reg state_4_4_13_lpi_3;
  reg state_4_4_50_lpi_3;
  reg state_4_4_12_lpi_3;
  reg state_4_4_51_lpi_3;
  reg state_4_4_11_lpi_3;
  reg state_4_4_52_lpi_3;
  reg state_4_4_10_lpi_3;
  reg state_4_4_53_lpi_3;
  reg state_4_4_9_lpi_3;
  reg state_4_4_54_lpi_3;
  reg state_4_4_8_lpi_3;
  reg state_4_4_55_lpi_3;
  reg state_4_4_7_lpi_3;
  reg state_4_4_56_lpi_3;
  reg state_4_4_6_lpi_3;
  reg state_4_4_57_lpi_3;
  reg state_4_4_5_lpi_3;
  reg state_4_4_58_lpi_3;
  reg state_4_4_4_lpi_3;
  reg state_4_4_59_lpi_3;
  reg state_4_4_3_lpi_3;
  reg state_4_4_60_lpi_3;
  reg state_4_4_2_lpi_3;
  reg state_4_4_61_lpi_3;
  reg state_4_4_1_lpi_3;
  reg state_4_4_62_lpi_3;
  reg state_4_4_0_lpi_3;
  reg state_4_4_63_lpi_3;
  reg [2:0] AD_P6_j_2_0_sva;
  reg state_0_31_lpi_6;
  reg state_0_32_lpi_6;
  reg state_0_30_lpi_6;
  reg state_0_33_lpi_6;
  reg state_0_29_lpi_6;
  reg state_0_34_lpi_6;
  reg state_0_28_lpi_6;
  reg state_0_35_lpi_6;
  reg state_0_27_lpi_6;
  reg state_0_36_lpi_6;
  reg state_0_26_lpi_6;
  reg state_0_37_lpi_6;
  reg state_0_25_lpi_6;
  reg state_0_38_lpi_6;
  reg state_0_24_lpi_6;
  reg state_0_39_lpi_6;
  reg state_0_23_lpi_6;
  reg state_0_40_lpi_6;
  reg state_0_22_lpi_6;
  reg state_0_41_lpi_6;
  reg state_0_21_lpi_6;
  reg state_0_42_lpi_6;
  reg state_0_20_lpi_6;
  reg state_0_43_lpi_6;
  reg state_0_19_lpi_6;
  reg state_0_44_lpi_6;
  reg state_0_18_lpi_6;
  reg state_0_45_lpi_6;
  reg state_0_17_lpi_6;
  reg state_0_46_lpi_6;
  reg state_0_16_lpi_6;
  reg state_0_47_lpi_6;
  reg state_0_15_lpi_6;
  reg state_0_48_lpi_6;
  reg state_0_14_lpi_6;
  reg state_0_49_lpi_6;
  reg state_0_13_lpi_6;
  reg state_0_50_lpi_6;
  reg state_0_12_lpi_6;
  reg state_0_51_lpi_6;
  reg state_0_11_lpi_6;
  reg state_0_52_lpi_6;
  reg state_0_10_lpi_6;
  reg state_0_53_lpi_6;
  reg state_0_9_lpi_6;
  reg state_0_54_lpi_6;
  reg state_0_8_lpi_6;
  reg state_0_55_lpi_6;
  reg state_0_7_lpi_6;
  reg state_0_56_lpi_6;
  reg state_0_6_lpi_6;
  reg state_0_57_lpi_6;
  reg state_0_5_lpi_6;
  reg state_0_58_lpi_6;
  reg state_0_4_lpi_6;
  reg state_0_59_lpi_6;
  reg state_0_3_lpi_6;
  reg state_0_60_lpi_6;
  reg state_0_2_lpi_6;
  reg state_0_61_lpi_6;
  reg state_0_1_lpi_6;
  reg state_0_62_lpi_6;
  reg state_0_0_lpi_6;
  reg state_0_63_lpi_6;
  reg state_2_0_1_lpi_6;
  reg state_2_1_1_lpi_6;
  reg state_2_2_1_lpi_6;
  reg state_2_3_1_lpi_6;
  reg state_2_4_1_lpi_6;
  reg state_2_5_1_lpi_6;
  reg state_2_6_1_lpi_6;
  reg state_2_7_1_lpi_6;
  reg state_1_1_31_0_lpi_4_31;
  reg state_1_1_31_0_lpi_4_30;
  reg state_1_1_31_0_lpi_4_29;
  reg state_1_1_31_0_lpi_4_28;
  reg state_1_1_31_0_lpi_4_27;
  reg state_1_1_31_0_lpi_4_26;
  reg state_1_1_31_0_lpi_4_25;
  reg state_1_1_31_0_lpi_4_24;
  reg state_1_1_31_0_lpi_4_23;
  reg state_1_1_31_0_lpi_4_22;
  reg state_1_1_31_0_lpi_4_21;
  reg state_1_1_31_0_lpi_4_20;
  reg state_1_1_31_0_lpi_4_19;
  reg state_1_1_31_0_lpi_4_18;
  reg state_1_1_31_0_lpi_4_17;
  reg state_1_1_31_0_lpi_4_16;
  reg state_1_1_31_0_lpi_4_15;
  reg state_1_1_31_0_lpi_4_14;
  reg state_1_1_31_0_lpi_4_13;
  reg state_1_1_31_0_lpi_4_12;
  reg state_1_1_31_0_lpi_4_11;
  reg state_1_1_31_0_lpi_4_10;
  reg state_1_1_31_0_lpi_4_9;
  reg state_1_1_31_0_lpi_4_8;
  reg state_1_1_31_0_lpi_4_7;
  reg state_1_1_31_0_lpi_4_6;
  reg state_1_1_31_0_lpi_4_5;
  reg state_1_1_31_0_lpi_4_4;
  reg state_1_1_31_0_lpi_4_3;
  reg state_1_1_31_0_lpi_4_2;
  reg state_1_1_31_0_lpi_4_1;
  reg state_1_1_31_0_lpi_4_0;
  reg state_1_1_63_32_lpi_4_31;
  reg state_1_1_63_32_lpi_4_30;
  reg state_1_1_63_32_lpi_4_29;
  reg state_1_1_63_32_lpi_4_28;
  reg state_1_1_63_32_lpi_4_27;
  reg state_1_1_63_32_lpi_4_26;
  reg state_1_1_63_32_lpi_4_25;
  reg state_1_1_63_32_lpi_4_24;
  reg state_1_1_63_32_lpi_4_23;
  reg state_1_1_63_32_lpi_4_22;
  reg state_1_1_63_32_lpi_4_21;
  reg state_1_1_63_32_lpi_4_20;
  reg state_1_1_63_32_lpi_4_19;
  reg state_1_1_63_32_lpi_4_18;
  reg state_1_1_63_32_lpi_4_17;
  reg state_1_1_63_32_lpi_4_16;
  reg state_1_1_63_32_lpi_4_15;
  reg state_1_1_63_32_lpi_4_14;
  reg state_1_1_63_32_lpi_4_13;
  reg state_1_1_63_32_lpi_4_12;
  reg state_1_1_63_32_lpi_4_11;
  reg state_1_1_63_32_lpi_4_10;
  reg state_1_1_63_32_lpi_4_9;
  reg state_1_1_63_32_lpi_4_8;
  reg state_1_1_63_32_lpi_4_7;
  reg state_1_1_63_32_lpi_4_6;
  reg state_1_1_63_32_lpi_4_5;
  reg state_1_1_63_32_lpi_4_4;
  reg state_1_1_63_32_lpi_4_3;
  reg state_1_1_63_32_lpi_4_2;
  reg state_1_1_63_32_lpi_4_1;
  reg state_1_1_63_32_lpi_4_0;
  wire ADLEN_ADLEN_xor_2_itm_mx0w0;
  wire state_0_0_sva_2_mx0w1;
  wire ciphertext_32_sva_mx0w2;
  wire data_out_rsci_idat_0_mx0w6;
  wire data_out_rsci_idat_0_mx0w7;
  wire ADLEN_ADLEN_xor_4_itm_mx0w0;
  wire state_0_1_sva_2_mx0w1;
  wire ciphertext_33_sva_mx0w2;
  wire data_out_rsci_idat_1_mx0w6;
  wire data_out_rsci_idat_1_mx0w7;
  wire ADLEN_ADLEN_xor_6_itm_mx0w0;
  wire state_0_2_sva_2_mx0w1;
  wire ciphertext_34_sva_mx0w2;
  wire data_out_rsci_idat_2_mx0w6;
  wire ADLEN_ADLEN_xor_8_itm_mx0w0;
  wire state_0_3_sva_2_mx0w1;
  wire ciphertext_35_sva_mx0w2;
  wire data_out_rsci_idat_3_mx0w6;
  wire ADLEN_ADLEN_xor_10_itm_mx0w0;
  wire state_0_4_sva_2_mx0w1;
  wire ciphertext_36_sva_mx0w2;
  wire data_out_rsci_idat_4_mx0w6;
  wire ADLEN_ADLEN_xor_12_itm_mx0w0;
  wire state_0_5_sva_2_mx0w1;
  wire ciphertext_37_sva_mx0w2;
  wire data_out_rsci_idat_5_mx0w6;
  wire ADLEN_ADLEN_xor_14_itm_mx0w0;
  wire state_0_6_sva_2_mx0w1;
  wire ciphertext_38_sva_mx0w2;
  wire data_out_rsci_idat_6_mx0w6;
  wire ADLEN_ADLEN_xor_16_itm_mx0w0;
  wire state_0_7_sva_2_mx0w1;
  wire ciphertext_39_sva_mx0w2;
  wire data_out_rsci_idat_7_mx0w6;
  wire ADLEN_ADLEN_xor_18_itm_mx0w0;
  wire state_0_8_sva_2_mx0w1;
  wire ciphertext_40_sva_mx0w2;
  wire data_out_rsci_idat_8_mx0w6;
  wire data_out_rsci_idat_8_mx0w7;
  wire ADLEN_ADLEN_xor_20_itm_mx0w0;
  wire state_0_9_sva_2_mx0w1;
  wire ciphertext_41_sva_mx0w2;
  wire data_out_rsci_idat_9_mx0w6;
  wire data_out_rsci_idat_9_mx0w7;
  wire ADLEN_ADLEN_xor_22_itm_mx0w0;
  wire state_0_10_sva_2_mx0w1;
  wire ciphertext_42_sva_mx0w2;
  wire data_out_rsci_idat_10_mx0w6;
  wire ADLEN_ADLEN_xor_24_itm_mx0w0;
  wire state_0_11_sva_2_mx0w1;
  wire ciphertext_43_sva_mx0w2;
  wire data_out_rsci_idat_11_mx0w6;
  wire ADLEN_ADLEN_xor_26_itm_mx0w0;
  wire state_0_12_sva_2_mx0w1;
  wire ciphertext_44_sva_mx0w2;
  wire data_out_rsci_idat_12_mx0w6;
  wire ADLEN_ADLEN_xor_28_itm_mx0w0;
  wire state_0_13_sva_2_mx0w1;
  wire ciphertext_45_sva_mx0w2;
  wire data_out_rsci_idat_13_mx0w6;
  wire ADLEN_ADLEN_xor_30_itm_mx0w0;
  wire state_0_14_sva_2_mx0w1;
  wire ciphertext_46_sva_mx0w2;
  wire data_out_rsci_idat_14_mx0w6;
  wire ADLEN_ADLEN_xor_32_itm_mx0w0;
  wire state_0_15_sva_2_mx0w1;
  wire ciphertext_47_sva_mx0w2;
  wire data_out_rsci_idat_15_mx0w6;
  wire ADLEN_ADLEN_xor_34_itm_mx0w0;
  wire state_0_16_sva_2_mx0w1;
  wire ciphertext_48_sva_mx0w2;
  wire data_out_rsci_idat_16_mx0w6;
  wire ADLEN_ADLEN_xor_36_itm_mx0w0;
  wire state_0_17_sva_2_mx0w1;
  wire ciphertext_49_sva_mx0w2;
  wire data_out_rsci_idat_17_mx0w6;
  wire ADLEN_ADLEN_xor_38_itm_mx0w0;
  wire state_0_18_sva_2_mx0w1;
  wire ciphertext_50_sva_mx0w2;
  wire data_out_rsci_idat_18_mx0w6;
  wire ADLEN_ADLEN_xor_40_itm_mx0w0;
  wire state_0_19_sva_2_mx0w1;
  wire ciphertext_51_sva_mx0w2;
  wire data_out_rsci_idat_19_mx0w6;
  wire ADLEN_ADLEN_xor_42_itm_mx0w0;
  wire state_0_20_sva_2_mx0w1;
  wire ciphertext_52_sva_mx0w2;
  wire data_out_rsci_idat_20_mx0w6;
  wire ADLEN_ADLEN_xor_44_itm_mx0w0;
  wire state_0_21_sva_2_mx0w1;
  wire ciphertext_53_sva_mx0w2;
  wire data_out_rsci_idat_21_mx0w6;
  wire ADLEN_ADLEN_xor_46_itm_mx0w0;
  wire state_0_22_sva_2_mx0w1;
  wire ciphertext_54_sva_mx0w2;
  wire data_out_rsci_idat_22_mx0w6;
  wire ADLEN_ADLEN_xor_48_itm_mx0w0;
  wire state_0_23_sva_2_mx0w1;
  wire ciphertext_55_sva_mx0w2;
  wire data_out_rsci_idat_23_mx0w6;
  wire ADLEN_ADLEN_xor_50_itm_mx0w0;
  wire state_0_24_sva_2_mx0w1;
  wire ciphertext_56_sva_mx0w2;
  wire data_out_rsci_idat_24_mx0w6;
  wire ADLEN_ADLEN_xor_52_itm_mx0w0;
  wire state_0_25_sva_2_mx0w1;
  wire ciphertext_57_sva_mx0w2;
  wire data_out_rsci_idat_25_mx0w6;
  wire ADLEN_ADLEN_xor_54_itm_mx0w0;
  wire state_0_26_sva_2_mx0w1;
  wire ciphertext_58_sva_mx0w2;
  wire ADLEN_ADLEN_xor_56_itm_mx0w0;
  wire state_0_27_sva_2_mx0w1;
  wire ciphertext_59_sva_mx0w2;
  wire ADLEN_ADLEN_xor_58_itm_mx0w0;
  wire state_0_28_sva_2_mx0w1;
  wire ciphertext_60_sva_mx0w2;
  wire ADLEN_ADLEN_xor_60_itm_mx0w0;
  wire state_0_29_sva_2_mx0w1;
  wire ciphertext_61_sva_mx0w2;
  wire ADLEN_ADLEN_xor_62_itm_mx0w0;
  wire state_0_30_sva_2_mx0w1;
  wire ciphertext_62_sva_mx0w2;
  wire ADLEN_ADLEN_xor_64_itm_mx0w0;
  wire state_0_31_sva_2_mx0w1;
  wire ciphertext_63_sva_mx0w2;
  wire state_0_4_sva_4_mx0w4;
  wire state_0_5_sva_4_mx0w4;
  wire state_0_6_sva_4_mx0w4;
  wire state_0_7_sva_4_mx0w4;
  wire state_4_16_sva_2_mx0w4;
  wire state_4_17_sva_2_mx0w4;
  wire state_4_18_sva_2_mx0w4;
  wire state_4_19_sva_2_mx0w4;
  wire state_4_2_sva_2_mx0w4;
  wire state_4_20_sva_2_mx0w4;
  wire state_4_21_sva_2_mx0w4;
  wire state_4_22_sva_2_mx0w4;
  wire state_4_4_23_sva_1_mx0w4;
  wire state_4_4_24_sva_1_mx0w4;
  wire state_4_25_sva_2_mx0w4;
  wire state_4_26_sva_2_mx0w4;
  wire state_4_27_sva_2_mx0w4;
  wire state_4_28_sva_2_mx0w4;
  wire state_4_29_sva_2_mx0w4;
  wire state_4_3_sva_2_mx0w4;
  wire state_4_30_sva_2_mx0w5;
  wire state_4_31_sva_2_mx0w5;
  wire state_4_4_sva_2_mx0w5;
  wire state_4_5_sva_2_mx0w5;
  wire state_4_6_sva_2_mx0w5;
  wire state_4_7_sva_2_mx0w5;
  wire state_4_32_sva_2_mx0w5;
  wire state_4_33_sva_2_mx0w5;
  wire state_4_34_sva_2_mx0w5;
  wire state_4_35_sva_2_mx0w5;
  wire state_4_36_sva_2_mx0w5;
  wire state_4_37_sva_2_mx0w5;
  wire state_4_38_sva_2_mx0w5;
  wire state_4_39_sva_2_mx0w5;
  wire state_4_40_sva_2_mx0w5;
  wire state_4_41_sva_2_mx0w5;
  wire state_4_42_sva_2_mx0w5;
  wire state_4_43_sva_2_mx0w5;
  wire state_4_44_sva_2_mx0w5;
  wire state_4_45_sva_2_mx0w5;
  wire state_4_46_sva_2_mx0w5;
  wire state_4_47_sva_2_mx0w5;
  wire state_4_48_sva_2_mx0w5;
  wire state_4_49_sva_2_mx0w5;
  wire state_4_50_sva_2_mx0w5;
  wire state_4_51_sva_2_mx0w5;
  wire state_4_52_sva_2_mx0w5;
  wire state_4_53_sva_2_mx0w5;
  wire state_4_54_sva_2_mx0w5;
  wire state_4_55_sva_2_mx0w5;
  wire state_4_56_sva_2_mx0w5;
  wire state_4_57_sva_2_mx0w5;
  wire state_4_8_sva_2_mx0w5;
  wire state_4_9_sva_2_mx0w5;
  wire state_0_8_sva_3_mx0w5;
  wire state_0_9_sva_3_mx0w5;
  wire state_3_0_sva_3_mx0w6;
  wire state_2_0_1_sva_4;
  wire state_3_1_sva_3_mx0w6;
  wire state_2_1_1_sva_4;
  wire state_3_10_sva_2_mx0w6;
  wire state_2_2_1_sva_4;
  wire state_3_11_sva_2_mx0w6;
  wire state_2_3_1_sva_4;
  wire state_3_12_sva_2_mx0w6;
  wire state_2_4_1_sva_4;
  wire state_3_13_sva_2_mx0w6;
  wire state_2_5_1_sva_4;
  wire state_3_14_sva_2_mx0w6;
  wire state_2_6_1_sva_4;
  wire state_3_15_sva_3_mx0w6;
  wire state_2_7_1_sva_4;
  wire ADLEN_i_7_0_sva_6_0_mx0c3;
  wire state_1_1_31_0_sva_1_31_1;
  wire state_1_1_31_0_sva_1_0_1;
  wire state_1_1_31_0_sva_1_30_1;
  wire state_1_1_31_0_sva_1_1_1;
  wire state_1_1_31_0_sva_1_29_1;
  wire state_1_1_31_0_sva_1_2_1;
  wire state_1_1_31_0_sva_1_28_1;
  wire state_1_1_31_0_sva_1_3_1;
  wire state_1_1_31_0_sva_1_27_1;
  wire state_1_1_31_0_sva_1_4_1;
  wire state_1_1_31_0_sva_1_26_1;
  wire state_1_1_31_0_sva_1_5_1;
  wire state_1_1_31_0_sva_1_25_1;
  wire state_1_1_31_0_sva_1_6_1;
  wire state_1_1_31_0_sva_1_24_1;
  wire state_1_1_31_0_sva_1_7_1;
  wire state_1_1_31_0_sva_1_23_1;
  wire state_1_1_31_0_sva_1_8_1;
  wire state_1_1_31_0_sva_1_22_1;
  wire state_1_1_31_0_sva_1_9_1;
  wire state_1_1_31_0_sva_1_21_1;
  wire state_1_1_31_0_sva_1_10_1;
  wire state_1_1_31_0_sva_1_20_1;
  wire state_1_1_31_0_sva_1_11_1;
  wire state_1_1_31_0_sva_1_19_1;
  wire state_1_1_31_0_sva_1_12_1;
  wire state_1_1_31_0_sva_1_18_1;
  wire state_1_1_31_0_sva_1_13_1;
  wire state_1_1_31_0_sva_1_17_1;
  wire state_1_1_31_0_sva_1_14_1;
  wire state_1_1_31_0_sva_1_16_1;
  wire state_1_1_31_0_sva_1_15_1;
  wire state_1_1_63_32_sva_1_31_1;
  wire state_1_1_63_32_sva_1_0_1;
  wire state_1_1_63_32_sva_1_30_1;
  wire state_1_1_63_32_sva_1_1_1;
  wire state_1_1_63_32_sva_1_29_1;
  wire state_1_1_63_32_sva_1_2_1;
  wire state_1_1_63_32_sva_1_28_1;
  wire state_1_1_63_32_sva_1_3_1;
  wire state_1_1_63_32_sva_1_27_1;
  wire state_1_1_63_32_sva_1_4_1;
  wire state_1_1_63_32_sva_1_26_1;
  wire state_1_1_63_32_sva_1_5_1;
  wire state_1_1_63_32_sva_1_25_1;
  wire state_1_1_63_32_sva_1_6_1;
  wire state_1_1_63_32_sva_1_24_1;
  wire state_1_1_63_32_sva_1_7_1;
  wire state_1_1_63_32_sva_1_23_1;
  wire state_1_1_63_32_sva_1_8_1;
  wire state_1_1_63_32_sva_1_22_1;
  wire state_1_1_63_32_sva_1_9_1;
  wire state_1_1_63_32_sva_1_21_1;
  wire state_1_1_63_32_sva_1_10_1;
  wire state_1_1_63_32_sva_1_20_1;
  wire state_1_1_63_32_sva_1_11_1;
  wire state_1_1_63_32_sva_1_19_1;
  wire state_1_1_63_32_sva_1_12_1;
  wire state_1_1_63_32_sva_1_18_1;
  wire state_1_1_63_32_sva_1_13_1;
  wire state_1_1_63_32_sva_1_17_1;
  wire state_1_1_63_32_sva_1_14_1;
  wire state_1_1_63_32_sva_1_16_1;
  wire state_1_1_63_32_sva_1_15_1;
  wire Encrypt_Top_sbox_and_2_cse_63_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_0_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_1_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_2_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_3_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_59_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_4_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_58_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_5_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_57_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_6_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_56_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_7_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_55_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_8_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_54_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_9_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_53_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_52_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_51_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_50_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_49_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_48_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_47_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_46_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_17_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_45_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_44_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_43_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_42_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_41_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_40_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_39_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_38_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_37_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_36_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_35_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_34_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_33_sva_1;
  wire Encrypt_Top_sbox_and_2_cse_32_sva_1;
  wire INIT_P12_INIT_P12_xor_8_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_7_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_6_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_5_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_4_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_3_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_2_psp_sva_1;
  wire INIT_P12_INIT_P12_xor_1_psp_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_63_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_0_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_62_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_1_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_61_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_2_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_60_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_3_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_59_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_4_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_58_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_5_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_57_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_6_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_56_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_7_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_55_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_8_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_54_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_9_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_53_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_10_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_52_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_11_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_51_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_12_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_50_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_13_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_49_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_14_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_48_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_15_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_47_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_16_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_46_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_17_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_45_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_18_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_44_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_19_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_43_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_20_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_42_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_21_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_41_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_22_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_40_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_23_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_39_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_24_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_38_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_25_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_37_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_26_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_36_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_27_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_35_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_28_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_34_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_29_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_33_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_30_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_32_sva_1;
  wire Encrypt_Top_sbox_and_1_cse_31_sva_1;
  wire state_3_16_sva_3_mx0w5;
  wire state_3_17_sva_3_mx0w5;
  wire state_3_27_sva_3_mx0w5;
  wire state_3_9_sva_3_mx0w5;
  wire state_4_60_sva_2_mx0w5;
  wire state_4_61_sva_2_mx0w5;
  wire state_4_62_sva_2_mx0w5;
  wire state_4_63_sva_2_mx0w5;
  wire state_3_18_sva_3_mx0w5;
  wire state_3_19_sva_3_mx0w4;
  wire state_3_2_sva_3_mx0w4;
  wire state_3_20_sva_3_mx0w4;
  wire state_3_21_sva_3_mx0w4;
  wire state_3_22_sva_3_mx0w4;
  wire state_3_23_sva_3_mx0w4;
  wire state_3_24_sva_3_mx0w4;
  wire state_3_25_sva_3_mx0w4;
  wire state_3_26_sva_3_mx0w4;
  wire state_3_28_sva_3_mx0w4;
  wire state_3_29_sva_3_mx0w4;
  wire state_3_3_sva_3_mx0w4;
  wire state_3_30_sva_3_mx0w4;
  wire state_3_31_sva_3_mx0w4;
  wire state_3_4_sva_3_mx0w5;
  wire state_3_5_sva_3_mx0w5;
  wire state_3_6_sva_3_mx0w5;
  wire state_3_7_sva_3_mx0w5;
  wire state_3_8_sva_3_mx0w5;
  wire state_4_58_sva_2_mx0w5;
  wire state_4_59_sva_2_mx0w5;
  wire state_4_0_sva_3;
  wire state_4_1_sva_3;
  wire state_4_10_sva_3;
  wire state_4_11_sva_3;
  wire state_4_12_sva_3;
  wire state_4_13_sva_3;
  wire state_4_14_sva_3;
  wire state_4_15_sva_3;
  wire [2:0] AD_P6_j_2_0_sva_2;
  wire [3:0] nl_AD_P6_j_2_0_sva_2;
  wire Encrypt_Top_sbox_1_and_cse_62_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_62_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_61_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_61_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_60_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_60_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_59_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_59_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_10_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_10_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_11_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_11_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_12_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_12_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_13_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_13_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_14_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_14_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_15_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_15_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_16_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_16_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_17_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_17_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_18_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_18_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_44_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_44_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_19_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_19_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_20_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_20_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_42_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_42_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_21_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_21_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_41_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_41_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_22_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_22_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_23_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_23_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_24_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_24_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_25_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_25_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_26_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_26_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_27_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_27_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_28_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_28_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_29_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_29_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_30_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_30_sva_1;
  wire Encrypt_Top_sbox_1_and_cse_31_sva_1;
  wire Encrypt_Top_sbox_2_and_2_cse_31_sva_1;
  wire AD_P6_AD_P6_xor_8_psp_sva_1;
  wire AD_P6_AD_P6_xor_7_psp_sva_1;
  wire AD_P6_AD_P6_xor_6_psp_sva_1;
  wire AD_P6_AD_P6_xor_5_psp_sva_1;
  wire AD_P6_AD_P6_xor_4_psp_sva_1;
  wire AD_P6_AD_P6_xor_3_psp_sva_1;
  wire AD_P6_AD_P6_xor_2_psp_sva_1;
  wire AD_P6_AD_P6_xor_1_psp_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_63_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_0_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_62_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_1_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_61_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_2_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_60_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_3_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_59_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_4_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_58_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_5_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_57_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_6_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_56_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_7_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_55_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_8_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_54_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_9_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_53_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_10_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_52_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_11_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_51_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_12_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_50_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_13_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_49_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_14_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_48_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_15_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_47_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_16_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_46_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_17_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_45_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_18_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_44_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_19_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_43_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_20_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_42_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_21_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_41_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_22_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_40_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_23_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_39_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_24_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_38_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_25_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_37_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_26_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_36_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_27_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_35_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_28_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_34_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_29_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_33_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_30_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_32_sva_1;
  wire Encrypt_Top_sbox_1_and_1_cse_31_sva_1;
  wire ENC_P6_ENC_P6_xor_8_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_7_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_6_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_5_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_4_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_3_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_2_psp_sva_1;
  wire ENC_P6_ENC_P6_xor_1_psp_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_0_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_1_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_2_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_3_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_4_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_5_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_6_sva_1;
  wire Encrypt_Top_sbox_2_and_1_cse_7_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_50_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_50_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_48_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_48_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_47_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_47_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_45_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_45_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_43_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_43_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_41_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_41_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_39_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_39_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_37_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_37_sva_1;
  wire Encrypt_Top_sbox_3_and_cse_36_sva_1;
  wire Encrypt_Top_sbox_3_and_2_cse_36_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_32_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_33_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_34_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_35_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_36_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_37_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_38_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_39_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_40_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_41_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_42_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_43_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_44_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_45_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_46_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_47_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_48_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_49_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_50_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_51_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_52_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_53_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_9_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_54_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_8_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_55_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_7_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_56_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_6_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_57_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_5_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_58_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_4_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_59_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_3_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_60_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_2_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_61_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_1_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_62_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_0_sva_1;
  wire Encrypt_Top_sbox_3_and_1_cse_63_sva_1;
  wire Encrypt_Top_sbox_2_and_516;
  wire Encrypt_Top_sbox_2_and_518;
  wire Encrypt_Top_sbox_1_and_516;
  wire Encrypt_Top_sbox_2_and_520;
  wire Encrypt_Top_sbox_2_and_522;
  wire Encrypt_Top_sbox_2_and_524;
  wire Encrypt_Top_sbox_2_and_526;
  wire Encrypt_Top_sbox_1_and_518;
  wire Encrypt_Top_sbox_2_and_528;
  wire Encrypt_Top_sbox_2_and_530;
  wire Encrypt_Top_sbox_2_and_532;
  wire Encrypt_Top_sbox_2_and_534;
  wire Encrypt_Top_sbox_1_and_520;
  wire Encrypt_Top_sbox_2_and_536;
  wire Encrypt_Top_sbox_2_and_538;
  wire Encrypt_Top_sbox_2_and_540;
  wire Encrypt_Top_sbox_2_and_542;
  wire Encrypt_Top_sbox_1_and_522;
  wire Encrypt_Top_sbox_2_and_544;
  wire Encrypt_Top_sbox_2_and_546;
  wire Encrypt_Top_sbox_2_and_548;
  wire Encrypt_Top_sbox_2_and_550;
  wire Encrypt_Top_sbox_1_and_524;
  wire Encrypt_Top_sbox_2_and_552;
  wire Encrypt_Top_sbox_2_and_554;
  wire Encrypt_Top_sbox_2_and_556;
  wire Encrypt_Top_sbox_2_and_558;
  wire Encrypt_Top_sbox_1_and_526;
  wire Encrypt_Top_sbox_2_and_560;
  wire Encrypt_Top_sbox_2_and_562;
  wire Encrypt_Top_sbox_2_and_564;
  wire Encrypt_Top_sbox_2_and_566;
  wire Encrypt_Top_sbox_1_and_528;
  wire Encrypt_Top_sbox_2_and_568;
  wire Encrypt_Top_sbox_2_and_570;
  wire Encrypt_Top_sbox_2_and_572;
  wire Encrypt_Top_sbox_2_and_574;
  wire Encrypt_Top_sbox_1_and_530;
  wire Encrypt_Top_sbox_2_and_576;
  wire Encrypt_Top_sbox_2_and_578;
  wire Encrypt_Top_sbox_2_and_580;
  wire Encrypt_Top_sbox_2_and_582;
  wire Encrypt_Top_sbox_1_and_532;
  wire Encrypt_Top_sbox_2_and_584;
  wire Encrypt_Top_sbox_2_and_586;
  wire Encrypt_Top_sbox_1_and_534;
  wire Encrypt_Top_sbox_2_and_588;
  wire Encrypt_Top_sbox_2_and_590;
  wire Encrypt_Top_sbox_1_and_536;
  wire Encrypt_Top_sbox_2_and_592;
  wire Encrypt_Top_sbox_2_and_594;
  wire Encrypt_Top_sbox_1_and_538;
  wire Encrypt_Top_sbox_2_and_596;
  wire Encrypt_Top_sbox_2_and_598;
  wire Encrypt_Top_sbox_1_and_540;
  wire Encrypt_Top_sbox_2_and_600;
  wire Encrypt_Top_sbox_2_and_602;
  wire Encrypt_Top_sbox_2_and_604;
  wire Encrypt_Top_sbox_2_and_606;
  wire Encrypt_Top_sbox_1_and_544;
  wire Encrypt_Top_sbox_2_and_608;
  wire Encrypt_Top_sbox_2_and_610;
  wire Encrypt_Top_sbox_2_and_612;
  wire Encrypt_Top_sbox_2_and_614;
  wire Encrypt_Top_sbox_1_and_548;
  wire Encrypt_Top_sbox_2_and_616;
  wire Encrypt_Top_sbox_2_and_618;
  wire Encrypt_Top_sbox_2_and_620;
  wire Encrypt_Top_sbox_2_and_622;
  wire Encrypt_Top_sbox_1_and_552;
  wire Encrypt_Top_sbox_2_and_624;
  wire Encrypt_Top_sbox_2_and_626;
  wire Encrypt_Top_sbox_2_and_628;
  wire Encrypt_Top_sbox_2_and_630;
  wire Encrypt_Top_sbox_1_and_556;
  wire Encrypt_Top_sbox_2_and_632;
  wire Encrypt_Top_sbox_2_and_634;
  wire Encrypt_Top_sbox_2_and_636;
  wire Encrypt_Top_sbox_2_and_638;
  wire Encrypt_Top_sbox_1_and_560;
  wire Encrypt_Top_sbox_2_and_640;
  wire Encrypt_Top_sbox_2_and_642;
  wire Encrypt_Top_sbox_2_and_644;
  wire Encrypt_Top_sbox_2_and_646;
  wire Encrypt_Top_sbox_1_and_564;
  wire Encrypt_Top_sbox_2_and_648;
  wire Encrypt_Top_sbox_2_and_650;
  wire Encrypt_Top_sbox_2_and_652;
  wire Encrypt_Top_sbox_2_and_654;
  wire Encrypt_Top_sbox_1_and_568;
  wire Encrypt_Top_sbox_2_and_656;
  wire Encrypt_Top_sbox_2_and_658;
  wire Encrypt_Top_sbox_2_and_660;
  wire Encrypt_Top_sbox_2_and_662;
  wire Encrypt_Top_sbox_1_and_572;
  wire Encrypt_Top_sbox_2_and_664;
  wire Encrypt_Top_sbox_2_and_666;
  wire Encrypt_Top_sbox_2_and_668;
  wire Encrypt_Top_sbox_2_and_670;
  wire Encrypt_Top_sbox_1_and_576;
  wire Encrypt_Top_sbox_2_and_672;
  wire Encrypt_Top_sbox_2_and_674;
  wire Encrypt_Top_sbox_2_and_676;
  wire Encrypt_Top_sbox_2_and_678;
  wire Encrypt_Top_sbox_1_and_580;
  wire Encrypt_Top_sbox_2_and_680;
  wire Encrypt_Top_sbox_2_and_682;
  wire Encrypt_Top_sbox_2_and_684;
  wire Encrypt_Top_sbox_2_and_686;
  wire Encrypt_Top_sbox_1_and_584;
  wire Encrypt_Top_sbox_2_and_688;
  wire Encrypt_Top_sbox_2_and_690;
  wire Encrypt_Top_sbox_2_and_692;
  wire Encrypt_Top_sbox_2_and_694;
  wire Encrypt_Top_sbox_1_and_588;
  wire Encrypt_Top_sbox_2_and_696;
  wire Encrypt_Top_sbox_2_and_698;
  wire Encrypt_Top_sbox_2_and_700;
  wire Encrypt_Top_sbox_2_and_702;
  wire Encrypt_Top_sbox_1_and_592;
  wire Encrypt_Top_sbox_2_and_704;
  wire Encrypt_Top_sbox_2_and_706;
  wire Encrypt_Top_sbox_2_and_708;
  wire Encrypt_Top_sbox_2_and_710;
  wire Encrypt_Top_sbox_1_and_596;
  wire Encrypt_Top_sbox_2_and_716;
  wire Encrypt_Top_sbox_2_and_718;
  wire Encrypt_Top_sbox_1_and_600;
  wire Encrypt_Top_sbox_2_and_724;
  wire Encrypt_Top_sbox_2_and_726;
  wire Encrypt_Top_sbox_1_and_604;
  wire Encrypt_Top_sbox_2_and_732;
  wire Encrypt_Top_sbox_2_and_734;
  wire Encrypt_Top_sbox_1_and_608;
  wire Encrypt_Top_sbox_2_and_740;
  wire Encrypt_Top_sbox_2_and_742;
  wire Encrypt_Top_sbox_1_and_612;
  wire Encrypt_Top_sbox_2_and_748;
  wire Encrypt_Top_sbox_2_and_750;
  wire Encrypt_Top_sbox_1_and_616;
  wire Encrypt_Top_sbox_2_and_752;
  wire Encrypt_Top_sbox_2_and_754;
  wire Encrypt_Top_sbox_2_and_756;
  wire Encrypt_Top_sbox_2_and_758;
  wire Encrypt_Top_sbox_1_and_620;
  wire Encrypt_Top_sbox_2_and_764;
  wire Encrypt_Top_sbox_2_and_766;
  wire Encrypt_Top_sbox_1_and_624;
  wire Encrypt_Top_sbox_1_and_628;
  wire Encrypt_Top_sbox_1_and_630;
  wire Encrypt_Top_sbox_1_and_632;
  wire Encrypt_Top_sbox_1_and_634;
  wire Encrypt_Top_sbox_1_and_636;
  wire Encrypt_Top_sbox_1_and_638;
  wire Encrypt_Top_sbox_1_and_640;
  wire Encrypt_Top_sbox_1_and_642;
  wire Encrypt_Top_sbox_1_and_652;
  wire Encrypt_Top_sbox_1_and_654;
  wire Encrypt_Top_sbox_1_and_656;
  wire Encrypt_Top_sbox_1_and_664;
  wire Encrypt_Top_sbox_1_and_666;
  wire Encrypt_Top_sbox_1_and_694;
  wire Encrypt_Top_sbox_1_and_728;
  wire Encrypt_Top_sbox_1_and_734;
  wire Encrypt_Top_sbox_1_and_756;
  wire Encrypt_Top_sbox_1_and_758;
  wire Encrypt_Top_sbox_1_and_760;
  wire Encrypt_Top_sbox_1_and_762;
  wire Encrypt_Top_sbox_1_and_764;
  wire Encrypt_Top_sbox_1_and_766;
  wire Encrypt_Top_sbox_1_and_768;
  wire Encrypt_Top_sbox_1_and_770;
  wire Encrypt_Top_sbox_1_and_784;
  wire Encrypt_Top_sbox_1_and_786;
  wire Encrypt_Top_sbox_1_and_788;
  wire Encrypt_Top_sbox_1_and_790;
  wire Encrypt_Top_sbox_1_and_792;
  wire Encrypt_Top_sbox_1_and_796;
  wire Encrypt_Top_sbox_1_and_798;
  wire Encrypt_Top_sbox_1_and_800;
  wire Encrypt_Top_sbox_1_and_802;
  wire Encrypt_Top_sbox_1_and_808;
  wire Encrypt_Top_sbox_1_and_816;
  wire Encrypt_Top_sbox_1_and_818;
  wire Encrypt_Top_sbox_1_and_820;
  wire Encrypt_Top_sbox_1_and_822;
  wire Encrypt_Top_sbox_1_and_824;
  wire Encrypt_Top_sbox_1_and_826;
  wire Encrypt_Top_sbox_1_and_828;
  wire Encrypt_Top_sbox_1_and_830;
  wire Encrypt_Top_sbox_1_and_832;
  wire Encrypt_Top_sbox_1_and_834;
  wire Encrypt_Top_sbox_1_and_836;
  wire Encrypt_Top_sbox_1_and_838;
  wire Encrypt_Top_sbox_1_and_840;
  wire Encrypt_Top_sbox_1_and_842;
  wire Encrypt_Top_sbox_1_and_844;
  wire Encrypt_Top_sbox_1_and_846;
  wire Encrypt_Top_sbox_1_and_848;
  wire Encrypt_Top_sbox_1_and_850;
  wire Encrypt_Top_sbox_1_and_852;
  wire Encrypt_Top_sbox_1_and_854;
  wire Encrypt_Top_sbox_1_and_856;
  wire Encrypt_Top_sbox_1_and_858;
  wire Encrypt_Top_sbox_1_and_860;
  wire Encrypt_Top_sbox_1_and_862;
  wire Encrypt_Top_sbox_1_and_864;
  wire Encrypt_Top_sbox_1_and_866;
  wire Encrypt_Top_sbox_1_and_868;
  wire Encrypt_Top_sbox_1_and_870;
  wire Encrypt_Top_sbox_1_and_872;
  wire Encrypt_Top_sbox_1_and_874;
  wire Encrypt_Top_sbox_1_and_876;
  wire Encrypt_Top_sbox_1_and_878;
  wire Encrypt_Top_sbox_1_and_880;
  wire Encrypt_Top_sbox_1_and_882;
  wire xor_cse;
  wire xor_cse_1;
  wire xor_cse_3;
  wire xor_cse_4;
  wire xor_cse_5;
  wire xor_cse_7;
  wire xor_cse_8;
  wire xor_cse_10;
  wire xor_cse_11;
  wire xor_cse_12;
  wire xor_cse_14;
  wire xor_cse_15;
  wire xor_cse_17;
  wire xor_cse_18;
  wire xor_cse_19;
  wire xor_cse_21;
  wire xor_cse_22;
  wire xor_cse_24;
  wire xor_cse_25;
  wire xor_cse_26;
  wire xor_cse_28;
  wire xor_cse_29;
  wire xor_cse_30;
  wire xor_cse_31;
  wire xor_cse_32;
  wire xor_cse_34;
  wire xor_cse_35;
  wire xor_cse_37;
  wire xor_cse_38;
  wire xor_cse_39;
  wire xor_cse_41;
  wire xor_cse_42;
  wire xor_cse_43;
  wire xor_cse_44;
  wire xor_cse_46;
  wire xor_cse_47;
  wire xor_cse_48;
  wire xor_cse_49;
  wire xor_cse_51;
  wire xor_cse_52;
  wire xor_cse_53;
  wire xor_cse_55;
  wire xor_cse_56;
  wire xor_cse_57;
  wire xor_cse_59;
  wire xor_cse_60;
  wire xor_cse_61;
  wire xor_cse_62;
  wire xor_cse_63;
  wire xor_cse_65;
  wire xor_cse_66;
  wire xor_cse_67;
  wire xor_cse_69;
  wire xor_cse_70;
  wire xor_cse_71;
  wire xor_cse_73;
  wire xor_cse_74;
  wire xor_cse_75;
  wire xor_cse_76;
  wire xor_cse_77;
  wire xor_cse_79;
  wire xor_cse_80;
  wire xor_cse_81;
  wire xor_cse_83;
  wire xor_cse_84;
  wire xor_cse_85;
  wire xor_cse_87;
  wire xor_cse_88;
  wire xor_cse_89;
  wire xor_cse_90;
  wire xor_cse_91;
  wire xor_cse_92;
  wire xor_cse_94;
  wire xor_cse_95;
  wire xor_cse_97;
  wire xor_cse_98;
  wire xor_cse_99;
  wire xor_cse_100;
  wire xor_cse_102;
  wire xor_cse_103;
  wire xor_cse_104;
  wire xor_cse_106;
  wire xor_cse_107;
  wire xor_cse_108;
  wire xor_cse_110;
  wire xor_cse_111;
  wire xor_cse_112;
  wire xor_cse_113;
  wire xor_cse_115;
  wire xor_cse_116;
  wire xor_cse_117;
  wire xor_cse_119;
  wire xor_cse_120;
  wire xor_cse_121;
  wire xor_cse_123;
  wire xor_cse_124;
  wire xor_cse_125;
  wire xor_cse_127;
  wire xor_cse_128;
  wire xor_cse_129;
  wire xor_cse_130;
  wire xor_cse_132;
  wire xor_cse_133;
  wire xor_cse_135;
  wire xor_cse_136;
  wire xor_cse_137;
  wire xor_cse_139;
  wire xor_cse_140;
  wire xor_cse_141;
  wire xor_cse_142;
  wire xor_cse_143;
  wire xor_cse_145;
  wire xor_cse_147;
  wire xor_cse_148;
  wire xor_cse_149;
  wire xor_cse_151;
  wire xor_cse_152;
  wire xor_cse_153;
  wire xor_cse_154;
  wire xor_cse_156;
  wire xor_cse_159;
  wire xor_cse_160;
  wire xor_cse_161;
  wire xor_cse_163;
  wire xor_cse_164;
  wire xor_cse_167;
  wire xor_cse_168;
  wire xor_cse_170;
  wire xor_cse_171;
  wire xor_cse_172;
  wire xor_cse_174;
  wire xor_cse_175;
  wire xor_cse_177;
  wire xor_cse_178;
  wire xor_cse_181;
  wire xor_cse_183;
  wire xor_cse_185;
  wire xor_cse_186;
  wire xor_cse_188;
  wire xor_cse_189;
  wire xor_cse_190;
  wire xor_cse_192;
  wire xor_cse_194;
  wire xor_cse_195;
  wire xor_cse_196;
  wire xor_cse_197;
  wire xor_cse_200;
  wire xor_cse_201;
  wire xor_cse_202;
  wire xor_cse_204;
  wire xor_cse_205;
  wire xor_cse_206;
  wire xor_cse_207;
  wire xor_cse_209;
  wire xor_cse_210;
  wire xor_cse_211;
  wire xor_cse_214;
  wire xor_cse_217;
  wire xor_cse_218;
  wire xor_cse_220;
  wire xor_cse_221;
  wire xor_cse_222;
  wire xor_cse_224;
  wire xor_cse_226;
  wire xor_cse_228;
  wire xor_cse_229;
  wire xor_cse_230;
  wire xor_cse_231;
  wire xor_cse_235;
  wire xor_cse_236;
  wire xor_cse_238;
  wire xor_cse_239;
  wire xor_cse_241;
  wire xor_cse_242;
  wire xor_cse_246;
  wire xor_cse_248;
  wire xor_cse_249;
  wire xor_cse_251;
  wire xor_cse_252;
  wire xor_cse_254;
  wire xor_cse_256;
  wire xor_cse_257;
  wire xor_cse_258;
  wire xor_cse_260;
  wire xor_cse_262;
  wire xor_cse_263;
  wire xor_cse_265;
  wire xor_cse_267;
  wire xor_cse_268;
  wire xor_cse_270;
  wire xor_cse_272;
  wire xor_cse_274;
  wire xor_cse_275;
  wire xor_cse_277;
  wire xor_cse_278;
  wire xor_cse_280;
  wire xor_cse_282;
  wire xor_cse_283;
  wire xor_cse_285;
  wire xor_cse_286;
  wire xor_cse_288;
  wire xor_cse_290;
  wire xor_cse_291;
  wire xor_cse_293;
  wire xor_cse_297;
  wire xor_cse_299;
  wire xor_cse_300;
  wire xor_cse_302;
  wire xor_cse_306;
  wire xor_cse_308;
  wire xor_cse_309;
  wire xor_cse_311;
  wire xor_cse_315;
  wire xor_cse_316;
  wire xor_cse_318;
  wire xor_cse_320;
  wire xor_cse_324;
  wire xor_cse_325;
  wire xor_cse_327;
  wire xor_cse_329;
  wire xor_cse_331;
  wire xor_cse_333;
  wire xor_cse_334;
  wire xor_cse_336;
  wire xor_cse_339;
  wire xor_cse_341;
  wire xor_cse_343;
  wire xor_cse_344;
  wire xor_cse_347;
  wire xor_cse_349;
  wire xor_cse_350;
  wire xor_cse_351;
  wire xor_cse_352;
  wire xor_cse_354;
  wire xor_cse_356;
  wire xor_cse_357;
  wire xor_cse_358;
  wire xor_cse_359;
  wire xor_cse_360;
  wire xor_cse_361;
  wire xor_cse_362;
  wire xor_cse_363;
  wire xor_cse_364;
  wire xor_cse_366;
  wire xor_cse_368;
  wire xor_cse_369;
  wire xor_cse_370;
  wire xor_cse_373;
  wire xor_cse_374;
  wire xor_cse_375;
  wire xor_cse_376;
  wire xor_cse_377;
  wire xor_cse_379;
  wire xor_cse_381;
  wire xor_cse_382;
  wire xor_cse_383;
  wire xor_cse_384;
  wire xor_cse_385;
  wire xor_cse_386;
  wire xor_cse_387;
  wire xor_cse_389;
  wire xor_cse_390;
  wire xor_cse_393;
  wire xor_cse_394;
  wire xor_cse_395;
  wire xor_cse_400;
  wire xor_cse_401;
  wire xor_cse_402;
  wire xor_cse_403;
  wire xor_cse_405;
  wire xor_cse_407;
  wire xor_cse_412;
  wire xor_cse_414;
  wire xor_cse_415;
  wire xor_cse_416;
  wire xor_cse_417;
  wire xor_cse_419;
  wire xor_cse_421;
  wire xor_cse_425;
  wire xor_cse_426;
  wire xor_cse_427;
  wire xor_cse_428;
  wire xor_cse_430;
  wire xor_cse_431;
  wire xor_cse_434;
  wire xor_cse_435;
  wire xor_cse_436;
  wire xor_cse_438;
  wire xor_cse_439;
  wire xor_cse_441;
  wire xor_cse_443;
  wire xor_cse_444;
  wire xor_cse_445;
  wire xor_cse_446;
  wire xor_cse_448;
  wire xor_cse_450;
  wire xor_cse_452;
  wire xor_cse_453;
  wire xor_cse_456;
  wire xor_cse_457;
  wire xor_cse_458;
  wire xor_cse_459;
  wire xor_cse_461;
  wire xor_cse_462;
  wire xor_cse_463;
  wire xor_cse_464;
  wire xor_cse_465;
  wire xor_cse_466;
  wire xor_cse_467;
  wire xor_cse_468;
  wire xor_cse_469;
  wire xor_cse_470;
  wire xor_cse_471;
  wire xor_cse_472;
  wire xor_cse_475;
  wire xor_cse_476;
  wire xor_cse_477;
  wire xor_cse_479;
  wire xor_cse_480;
  wire xor_cse_481;
  wire xor_cse_482;
  wire xor_cse_483;
  wire xor_cse_487;
  wire xor_cse_488;
  wire xor_cse_490;
  wire xor_cse_491;
  wire xor_cse_492;
  wire xor_cse_494;
  wire xor_cse_495;
  wire xor_cse_496;
  wire xor_cse_498;
  wire xor_cse_499;
  wire xor_cse_500;
  wire xor_cse_502;
  wire xor_cse_503;
  wire xor_cse_504;
  wire xor_cse_505;
  wire xor_cse_506;
  wire xor_cse_507;
  wire xor_cse_509;
  wire xor_cse_511;
  wire xor_cse_513;
  wire xor_cse_514;
  wire xor_cse_515;
  wire xor_cse_516;
  wire xor_cse_519;
  wire xor_cse_520;
  wire xor_cse_521;
  wire xor_cse_522;
  wire xor_cse_525;
  wire xor_cse_526;
  wire xor_cse_527;
  wire xor_cse_528;
  wire xor_cse_529;
  wire xor_cse_532;
  wire xor_cse_535;
  wire xor_cse_536;
  wire xor_cse_538;
  wire xor_cse_539;
  wire xor_cse_542;
  wire xor_cse_543;
  wire xor_cse_544;
  wire xor_cse_546;
  wire xor_cse_547;
  wire xor_cse_548;
  wire xor_cse_549;
  wire xor_cse_551;
  wire xor_cse_552;
  wire xor_cse_553;
  wire xor_cse_554;
  wire xor_cse_556;
  wire xor_cse_557;
  wire xor_cse_558;
  wire xor_cse_559;
  wire xor_cse_561;
  wire xor_cse_562;
  wire xor_cse_565;
  wire xor_cse_566;
  wire xor_cse_568;
  wire xor_cse_569;
  wire xor_cse_570;
  wire xor_cse_571;
  wire xor_cse_574;
  wire xor_cse_575;
  wire xor_cse_576;
  wire xor_cse_577;
  wire xor_cse_581;
  wire xor_cse_585;
  wire xor_cse_586;
  wire xor_cse_587;
  wire xor_cse_588;
  wire xor_cse_589;
  wire xor_cse_590;
  wire xor_cse_591;
  wire xor_cse_594;
  wire xor_cse_595;
  wire xor_cse_597;
  wire xor_cse_601;
  wire xor_cse_602;
  wire xor_cse_603;
  wire xor_cse_604;
  wire xor_cse_605;
  wire xor_cse_606;
  wire xor_cse_607;
  wire xor_cse_608;
  wire xor_cse_609;
  wire xor_cse_610;
  wire xor_cse_613;
  wire xor_cse_614;
  wire xor_cse_616;
  wire xor_cse_618;
  wire xor_cse_619;
  wire xor_cse_621;
  wire xor_cse_624;
  wire xor_cse_628;
  wire xor_cse_629;
  wire xor_cse_631;
  wire xor_cse_633;
  wire xor_cse_634;
  wire xor_cse_635;
  wire xor_cse_636;
  wire xor_cse_637;
  wire xor_cse_641;
  wire xor_cse_643;
  wire xor_cse_645;
  wire xor_cse_650;
  wire xor_cse_651;
  wire xor_cse_653;
  wire xor_cse_656;
  wire xor_cse_659;
  wire xor_cse_664;
  wire xor_cse_667;
  wire xor_cse_672;
  wire xor_cse_673;
  wire xor_cse_676;
  wire xor_cse_680;
  wire xor_cse_683;
  wire xor_cse_685;
  wire xor_cse_689;
  wire xor_cse_690;
  wire xor_cse_691;
  wire xor_cse_694;
  wire xor_cse_698;
  wire xor_cse_701;
  wire xor_cse_702;
  wire xor_cse_705;
  wire xor_cse_708;
  wire xor_cse_709;
  wire xor_cse_713;
  wire xor_cse_716;
  wire xor_cse_717;
  wire xor_cse_721;
  wire xor_cse_722;
  wire xor_cse_724;
  wire xor_cse_725;
  wire xor_cse_726;
  wire xor_cse_730;
  wire xor_cse_732;
  wire xor_cse_734;
  wire xor_cse_735;
  wire xor_cse_736;
  wire xor_cse_739;
  wire xor_cse_740;
  wire xor_cse_742;
  wire xor_cse_743;
  wire xor_cse_746;
  wire xor_cse_748;
  wire xor_cse_749;
  wire xor_cse_752;
  wire xor_cse_753;
  wire xor_cse_754;
  wire xor_cse_755;
  wire xor_cse_759;
  wire xor_cse_760;
  wire xor_cse_763;
  wire xor_cse_764;
  wire xor_cse_767;
  wire xor_cse_769;
  wire xor_cse_770;
  wire xor_cse_771;
  wire xor_cse_775;
  wire xor_cse_776;
  wire xor_cse_777;
  wire xor_cse_782;
  wire xor_cse_783;
  wire xor_cse_784;
  wire xor_cse_788;
  wire xor_cse_789;
  wire xor_cse_790;
  wire xor_cse_792;
  wire xor_cse_794;
  wire xor_cse_795;
  wire xor_cse_796;
  wire xor_cse_797;
  wire xor_cse_799;
  wire xor_cse_801;
  wire xor_cse_802;
  wire xor_cse_805;
  wire xor_cse_806;
  wire xor_cse_807;
  wire xor_cse_808;
  wire xor_cse_809;
  wire xor_cse_812;
  wire xor_cse_813;
  wire xor_cse_814;
  wire xor_cse_817;
  wire xor_cse_820;
  wire xor_cse_821;
  wire xor_cse_822;
  wire xor_cse_825;
  wire xor_cse_826;
  wire xor_cse_827;
  wire xor_cse_829;
  wire xor_cse_832;
  wire xor_cse_833;
  wire xor_cse_834;
  wire xor_cse_835;
  wire xor_cse_839;
  wire xor_cse_842;
  wire xor_cse_845;
  wire xor_cse_847;
  wire xor_cse_850;
  wire xor_cse_851;
  wire xor_cse_852;
  wire xor_cse_854;
  wire xor_cse_858;
  wire xor_cse_859;
  wire xor_cse_861;
  wire xor_cse_866;
  wire xor_cse_867;
  wire xor_cse_868;
  wire xor_cse_871;
  wire xor_cse_875;
  wire xor_cse_877;
  wire xor_cse_878;
  wire xor_cse_880;
  wire xor_cse_887;
  wire xor_cse_888;
  wire xor_cse_890;
  wire xor_cse_895;
  wire xor_cse_897;
  wire xor_cse_899;
  wire xor_cse_900;
  wire xor_cse_905;
  wire xor_cse_906;
  wire xor_cse_909;
  wire xor_cse_910;
  wire xor_cse_912;
  wire xor_cse_915;
  wire xor_cse_920;
  wire xor_cse_923;
  wire xor_cse_924;
  wire xor_cse_926;
  wire xor_cse_927;
  wire xor_cse_928;
  wire xor_cse_932;
  wire xor_cse_933;
  wire xor_cse_935;
  wire xor_cse_936;
  wire xor_cse_943;
  wire xor_cse_944;
  wire xor_cse_947;
  wire xor_cse_948;
  wire xor_cse_950;
  wire xor_cse_951;
  wire xor_cse_953;
  wire xor_cse_955;
  wire xor_cse_958;
  wire xor_cse_961;
  wire xor_cse_967;
  wire xor_cse_970;
  wire xor_cse_977;
  wire xor_cse_981;
  wire xor_cse_983;
  wire xor_cse_985;
  wire xor_cse_990;
  wire xor_cse_996;
  wire xor_cse_1000;
  wire xor_cse_1009;
  wire xor_cse_1016;
  wire xor_cse_1017;
  wire xor_cse_1018;
  wire xor_cse_1021;
  wire xor_cse_1030;
  wire xor_cse_1031;
  wire xor_cse_1034;
  wire xor_cse_1037;
  wire xor_cse_1041;
  wire xor_cse_1046;
  wire xor_cse_1050;
  wire xor_cse_1055;
  wire xor_cse_1059;
  wire xor_cse_1064;
  wire xor_cse_1068;
  wire xor_cse_1077;
  wire xor_cse_1078;
  wire xor_cse_1085;
  wire xor_cse_1086;
  wire xor_cse_1087;
  wire xor_cse_1095;
  wire xor_cse_1096;
  wire xor_cse_1097;
  wire xor_cse_1103;
  wire xor_cse_1108;
  wire xor_cse_1134;
  wire xor_cse_1144;
  wire xor_cse_1161;
  wire xor_cse_1162;
  wire xor_cse_1167;
  wire xor_cse_1171;
  wire xor_cse_1172;
  wire xor_cse_1187;
  wire xor_cse_1188;
  wire xor_cse_1193;
  wire xor_cse_1293;
  wire xor_cse_1299;
  wire xor_cse_1300;
  wire xor_cse_1301;
  wire xor_cse_1303;
  wire xor_cse_1306;
  wire xor_cse_1309;
  wire xor_cse_1310;
  wire xor_cse_1311;
  wire xor_cse_1317;
  wire xor_cse_1324;
  wire xor_cse_1325;
  wire xor_cse_1332;
  wire xor_cse_1341;
  wire xor_cse_1350;
  wire xor_cse_1351;
  wire xor_cse_1357;
  wire xor_cse_1358;
  wire xor_cse_1360;
  wire xor_cse_1361;
  wire xor_cse_1363;
  wire xor_cse_1364;
  wire xor_cse_1366;
  wire xor_cse_1367;
  wire xor_cse_1368;
  wire xor_cse_1371;
  wire xor_cse_1374;
  wire xor_cse_1375;
  wire xor_cse_1378;
  wire xor_cse_1381;
  wire xor_cse_1382;
  wire xor_cse_1384;
  wire xor_cse_1385;
  wire xor_cse_1386;
  wire xor_cse_1388;
  wire xor_cse_1389;
  wire xor_cse_1391;
  wire xor_cse_1392;
  wire xor_cse_1393;
  wire xor_cse_1396;
  wire xor_cse_1399;
  wire xor_cse_1400;
  wire xor_cse_1403;
  wire xor_cse_1406;
  wire xor_cse_1408;
  wire xor_cse_1409;
  wire xor_cse_1410;
  wire xor_cse_1412;
  wire xor_cse_1413;
  wire xor_cse_1415;
  wire xor_cse_1416;
  wire xor_cse_1417;
  wire xor_cse_1418;
  wire xor_cse_1419;
  wire xor_cse_1420;
  wire xor_cse_1423;
  wire xor_cse_1426;
  wire xor_cse_1429;
  wire xor_cse_1430;
  wire xor_cse_1431;
  wire xor_cse_1433;
  wire xor_cse_1434;
  wire xor_cse_1436;
  wire xor_cse_1437;
  wire xor_cse_1439;
  wire xor_cse_1441;
  wire xor_cse_1446;
  wire xor_cse_1451;
  wire xor_cse_1453;
  wire xor_cse_1454;
  wire xor_cse_1455;
  wire xor_cse_1456;
  wire xor_cse_1463;
  wire xor_cse_1465;
  wire xor_cse_1468;
  wire xor_cse_1475;
  wire xor_cse_1477;
  wire xor_cse_1478;
  wire xor_cse_1479;
  wire xor_cse_1482;
  wire xor_cse_1485;
  wire xor_cse_1487;
  wire xor_cse_1488;
  wire xor_cse_1489;
  wire xor_cse_1490;
  wire xor_cse_1491;
  wire xor_cse_1492;
  wire xor_cse_1497;
  wire xor_cse_1498;
  wire xor_cse_1499;
  wire xor_cse_1503;
  wire xor_cse_1505;
  wire xor_cse_1511;
  wire xor_cse_1512;
  wire xor_cse_1513;
  wire xor_cse_1514;
  wire xor_cse_1515;
  wire xor_cse_1517;
  wire xor_cse_1519;
  wire xor_cse_1525;
  wire xor_cse_1526;
  wire xor_cse_1527;
  wire xor_cse_1528;
  wire xor_cse_1531;
  wire xor_cse_1532;
  wire xor_cse_1533;
  wire xor_cse_1535;
  wire xor_cse_1538;
  wire xor_cse_1540;
  wire xor_cse_1541;
  wire xor_cse_1542;
  wire xor_cse_1543;
  wire xor_cse_1545;
  wire xor_cse_1546;
  wire xor_cse_1550;
  wire xor_cse_1551;
  wire xor_cse_1555;
  wire xor_cse_1556;
  wire xor_cse_1558;
  wire xor_cse_1559;
  wire xor_cse_1562;
  wire xor_cse_1564;
  wire xor_cse_1565;
  wire xor_cse_1566;
  wire xor_cse_1567;
  wire xor_cse_1568;
  wire xor_cse_1569;
  wire xor_cse_1571;
  wire xor_cse_1572;
  wire xor_cse_1574;
  wire xor_cse_1575;
  wire xor_cse_1576;
  wire xor_cse_1577;
  wire xor_cse_1578;
  wire xor_cse_1580;
  wire xor_cse_1581;
  wire xor_cse_1582;
  wire xor_cse_1583;
  wire xor_cse_1584;
  wire xor_cse_1585;
  wire xor_cse_1586;
  wire xor_cse_1587;
  wire xor_cse_1588;
  wire xor_cse_1589;
  wire xor_cse_1591;
  wire xor_cse_1595;
  wire xor_cse_1596;
  wire xor_cse_1598;
  wire xor_cse_1600;
  wire xor_cse_1601;
  wire xor_cse_1602;
  wire xor_cse_1604;
  wire xor_cse_1609;
  wire xor_cse_1614;
  wire xor_cse_1617;
  wire xor_cse_1623;
  wire xor_cse_1629;
  wire xor_cse_1637;
  wire xor_cse_1641;
  wire xor_cse_1642;
  wire xor_cse_1647;
  wire xor_cse_1648;
  wire xor_cse_1649;
  wire xor_cse_1650;
  wire xor_cse_1660;
  wire xor_cse_1662;
  wire xor_cse_1680;
  wire xor_cse_1690;
  wire xor_cse_1696;
  wire xor_cse_1702;
  wire xor_cse_1708;
  wire xor_cse_1714;
  wire xor_cse_1731;
  wire xor_cse_1732;
  wire xor_cse_1733;
  wire xor_cse_1734;
  wire xor_cse_1735;
  wire xor_cse_1736;
  wire xor_cse_1737;
  wire xor_cse_1738;
  wire xor_cse_1739;
  wire xor_cse_1740;
  wire xor_cse_1741;
  wire xor_cse_1742;
  wire xor_cse_1743;
  wire xor_cse_1744;
  wire xor_cse_1745;
  wire xor_cse_1746;
  wire xor_cse_1747;
  wire xor_cse_1748;
  wire xor_cse_1749;
  wire xor_cse_1750;
  wire xor_cse_1751;
  wire xor_cse_1752;
  wire xor_cse_1753;
  wire xor_cse_1754;
  wire xor_cse_1755;
  wire xor_cse_1756;
  wire xor_cse_1757;
  wire xor_cse_1758;
  wire xor_cse_1759;
  wire xor_cse_1760;
  wire xor_cse_1761;
  wire xor_cse_1762;
  wire xor_cse_1763;
  wire xor_cse_1764;
  wire xor_cse_1765;
  wire xor_cse_1766;
  wire xor_cse_1767;
  wire xor_cse_1768;
  wire xor_cse_1769;
  wire xor_cse_1770;
  wire xor_cse_1771;
  wire xor_cse_1772;
  wire xor_cse_1773;
  wire xor_cse_1774;
  wire xor_cse_1775;
  wire xor_cse_1776;
  wire xor_cse_1777;
  wire xor_cse_1778;
  wire xor_cse_1779;
  wire xor_cse_1780;
  wire xor_cse_1781;
  wire xor_cse_1782;
  wire xor_cse_1783;
  wire xor_cse_1784;
  wire xor_cse_1785;
  wire xor_cse_1786;
  wire xor_cse_1787;
  wire xor_cse_1788;
  wire xor_cse_1789;
  wire xor_cse_1790;
  wire xor_cse_1792;
  wire xor_cse_1793;
  wire xor_cse_1794;
  wire xor_cse_1795;
  wire xor_cse_1796;
  wire xor_cse_1797;
  wire xor_cse_1798;
  wire xor_cse_1799;
  wire xor_cse_1800;
  wire xor_cse_1801;
  wire xor_cse_1802;
  wire xor_cse_1803;
  wire xor_cse_1804;
  wire xor_cse_1835;
  wire xor_cse_1838;
  wire xor_cse_1842;
  wire xor_cse_1843;
  wire xor_cse_1844;
  wire xor_cse_1845;
  wire xor_cse_1849;
  wire xor_cse_1852;
  wire xor_cse_1853;
  wire xor_cse_1854;
  wire xor_cse_1855;
  wire xor_cse_1859;
  wire xor_cse_1860;
  wire xor_cse_1861;
  wire xor_cse_1862;
  wire xor_cse_1864;
  wire xor_cse_1865;
  wire xor_cse_1868;
  wire xor_cse_1871;
  wire xor_cse_1874;
  wire xor_cse_1877;
  wire xor_cse_1880;
  wire xor_cse_1881;
  wire xor_cse_1882;
  wire xor_cse_1883;
  wire xor_cse_1886;
  wire xor_cse_1889;
  wire xor_cse_1892;
  wire xor_cse_1895;
  wire xor_cse_1898;
  wire xor_cse_1899;
  wire xor_cse_1900;
  wire xor_cse_1901;
  wire xor_cse_1904;
  wire xor_cse_1907;
  wire xor_cse_1910;
  wire xor_cse_1913;
  wire xor_cse_1916;
  wire xor_cse_1919;
  wire xor_cse_1922;
  wire xor_cse_1925;
  wire xor_cse_1928;
  wire xor_cse_1931;
  wire xor_cse_1936;
  wire xor_cse_1941;
  wire xor_cse_1945;
  wire xor_cse_1946;
  wire xor_cse_1951;
  wire xor_cse_1955;
  wire xor_cse_1960;
  wire xor_cse_1963;
  wire xor_cse_1966;
  wire xor_cse_1969;
  wire xor_cse_1970;
  wire xor_cse_1973;
  wire xor_cse_1976;
  wire xor_cse_1979;
  wire xor_cse_1982;
  wire xor_cse_1985;
  wire xor_cse_1988;
  wire xor_cse_1991;
  wire xor_cse_1995;
  wire xor_cse_1996;
  wire xor_cse_1997;
  wire xor_cse_1998;
  wire xor_cse_2001;
  wire xor_cse_2005;
  wire xor_cse_2006;
  wire xor_cse_2007;
  wire xor_cse_2008;
  wire xor_cse_2013;
  wire xor_cse_2017;
  wire xor_cse_2018;
  wire xor_cse_2019;
  wire xor_cse_2021;
  wire xor_cse_2022;
  wire xor_cse_2024;
  wire xor_cse_2025;
  wire xor_cse_2029;
  wire xor_cse_2030;
  wire xor_cse_2032;
  wire xor_cse_2033;
  wire xor_cse_2036;
  wire xor_cse_2040;
  wire xor_cse_2041;
  wire xor_cse_2042;
  wire xor_cse_2044;
  wire xor_cse_2045;
  wire xor_cse_2046;
  wire xor_cse_2047;
  wire xor_cse_2053;
  wire xor_cse_2054;
  wire xor_cse_2055;
  wire xor_cse_2065;
  wire xor_cse_2069;
  wire xor_cse_2086;
  wire xor_cse_2089;
  wire xor_cse_2091;
  wire xor_cse_2095;
  wire xor_cse_2096;
  wire xor_cse_2098;
  wire xor_cse_2100;
  wire xor_cse_2104;
  wire xor_cse_2106;
  wire xor_cse_2108;
  wire xor_cse_2109;
  wire xor_cse_2110;
  wire xor_cse_2111;
  wire xor_cse_2112;
  wire xor_cse_2113;
  wire xor_cse_2114;
  wire xor_cse_2115;
  wire xor_cse_2118;
  wire xor_cse_2120;
  wire xor_cse_2123;
  wire xor_cse_2126;
  wire xor_cse_2129;
  wire xor_cse_2131;
  wire xor_cse_2132;
  wire xor_cse_2134;
  wire xor_cse_2137;
  wire xor_cse_2138;
  wire xor_cse_2142;
  wire xor_cse_2145;
  wire xor_cse_2148;
  wire xor_cse_2151;
  wire xor_cse_2153;
  wire xor_cse_2157;
  wire xor_cse_2159;
  wire xor_cse_2162;
  wire xor_cse_2167;
  wire xor_cse_2168;
  wire xor_cse_2172;
  wire xor_cse_2176;
  wire xor_cse_2178;
  wire xor_cse_2182;
  wire xor_cse_2184;
  wire xor_cse_2187;
  wire xor_cse_2190;
  wire xor_cse_2192;
  wire xor_cse_2196;
  wire xor_cse_2197;
  wire xor_cse_2201;
  wire xor_cse_2204;
  wire xor_cse_2205;
  wire xor_cse_2209;
  wire xor_cse_2213;
  wire xor_cse_2215;
  wire xor_cse_2219;
  wire xor_cse_2221;
  wire xor_cse_2224;
  wire xor_cse_2227;
  wire xor_cse_2229;
  wire xor_cse_2230;
  wire xor_cse_2234;
  wire xor_cse_2237;
  wire xor_cse_2241;
  wire xor_cse_2242;
  wire xor_cse_2243;
  wire xor_cse_2245;
  wire xor_cse_2249;
  wire xor_cse_2252;
  wire xor_cse_2255;
  wire xor_cse_2256;
  wire xor_cse_2258;
  wire xor_cse_2259;
  wire xor_cse_2261;
  wire xor_cse_2262;
  wire xor_cse_2264;
  wire xor_cse_2265;
  wire xor_cse_2268;
  wire xor_cse_2269;
  wire xor_cse_2271;
  wire xor_cse_2272;
  wire xor_cse_2274;
  wire xor_cse_2278;
  wire xor_cse_2279;
  wire xor_cse_2280;
  wire xor_cse_2281;
  wire xor_cse_2283;
  wire xor_cse_2286;
  wire xor_cse_2289;
  wire xor_cse_2290;
  wire xor_cse_2293;
  wire xor_cse_2297;
  wire xor_cse_2298;
  wire xor_cse_2299;
  wire xor_cse_2302;
  wire xor_cse_2308;
  wire xor_cse_2309;
  wire xor_cse_2313;
  wire xor_cse_2315;
  wire xor_cse_2316;
  wire xor_cse_2319;
  wire xor_cse_2321;
  wire xor_cse_2323;
  wire xor_cse_2327;
  wire xor_cse_2330;
  wire xor_cse_2331;
  wire xor_cse_2333;
  wire xor_cse_2336;
  wire xor_cse_2340;
  wire xor_cse_2342;
  wire xor_cse_2344;
  wire xor_cse_2351;
  wire xor_cse_2352;
  wire xor_cse_2356;
  wire xor_cse_2360;
  wire xor_cse_2361;
  wire xor_cse_2366;
  wire xor_cse_2367;
  wire xor_cse_2370;
  wire xor_cse_2371;
  wire xor_cse_2372;
  wire xor_cse_2373;
  wire xor_cse_2374;
  wire xor_cse_2375;
  wire xor_cse_2379;
  wire xor_cse_2383;
  wire xor_cse_2387;
  wire xor_cse_2388;
  wire xor_cse_2389;
  wire xor_cse_2390;
  wire xor_cse_2393;
  wire xor_cse_2395;
  wire xor_cse_2396;
  wire xor_cse_2397;
  wire xor_cse_2398;
  wire xor_cse_2399;
  wire xor_cse_2400;
  wire xor_cse_2405;
  wire xor_cse_2406;
  wire xor_cse_2407;
  wire xor_cse_2408;
  wire xor_cse_2413;
  wire xor_cse_2414;
  wire xor_cse_2416;
  wire xor_cse_2421;
  wire xor_cse_2422;
  wire xor_cse_2423;
  wire xor_cse_2426;
  wire xor_cse_2427;
  wire xor_cse_2429;
  wire xor_cse_2435;
  wire xor_cse_2436;
  wire xor_cse_2439;
  wire xor_cse_2442;
  wire xor_cse_2443;
  wire xor_cse_2448;
  wire xor_cse_2452;
  wire xor_cse_2457;
  wire xor_cse_2461;
  wire xor_cse_2463;
  wire xor_cse_2468;
  wire xor_cse_2469;
  wire xor_cse_2472;
  wire xor_cse_2476;
  wire xor_cse_2477;
  wire xor_cse_2488;
  wire xor_cse_2505;
  wire xor_cse_2510;
  wire xor_cse_2516;
  wire xor_cse_2543;
  wire xor_cse_2544;
  wire xor_cse_2545;
  wire xor_cse_2549;
  wire xor_cse_2559;
  wire xor_cse_2565;
  wire xor_cse_2598;
  wire xor_cse_2602;
  wire xor_cse_2604;
  wire xor_cse_2608;
  wire xor_cse_2610;
  wire xor_cse_2612;
  wire xor_cse_2618;
  wire xor_cse_2620;
  wire xor_cse_2625;
  wire xor_cse_2626;
  wire xor_cse_2629;
  wire xor_cse_2641;
  wire xor_cse_2688;
  wire xor_cse_2707;
  wire xor_cse_2771;
  wire xor_cse_2791;
  wire xor_cse_2799;
  wire xor_cse_2808;
  wire xor_cse_2814;
  wire xor_cse_2822;
  wire xor_cse_2827;
  wire xor_cse_2830;
  wire xor_cse_2836;
  wire xor_cse_2848;
  wire xor_cse_2855;
  wire xor_cse_2868;
  wire xor_cse_2887;
  wire xor_cse_2889;
  wire xor_cse_2891;
  wire xor_cse_2893;
  wire xor_cse_2895;
  wire xor_cse_2897;
  wire xor_cse_2903;
  wire xor_cse_2906;
  wire xor_cse_2909;
  wire xor_cse_2912;
  reg [2:0] ADLEN_i_7_0_sva_6_4;
  reg [3:0] ADLEN_i_7_0_sva_3_0;
  wire [7:0] ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1;
  wire [7:0] ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1;
  reg state_3_3_31_0_sva_31;
  reg state_3_3_31_0_sva_30;
  reg state_3_3_31_0_sva_29;
  reg state_3_3_31_0_sva_28;
  reg state_3_3_31_0_sva_27;
  reg state_3_3_31_0_sva_26;
  reg state_3_3_31_0_sva_25;
  reg state_3_3_31_0_sva_24;
  reg state_3_3_31_0_sva_23;
  reg state_3_3_31_0_sva_22;
  reg state_3_3_31_0_sva_21;
  reg state_3_3_31_0_sva_20;
  reg state_3_3_31_0_sva_19;
  reg state_3_3_31_0_sva_18;
  reg state_3_3_31_0_sva_17;
  reg state_3_3_31_0_sva_16;
  reg state_3_3_31_0_sva_15;
  reg state_3_3_31_0_sva_14;
  reg state_3_3_31_0_sva_13;
  reg state_3_3_31_0_sva_12;
  reg state_3_3_31_0_sva_11;
  reg state_3_3_31_0_sva_10;
  reg state_3_3_31_0_sva_9;
  reg state_3_3_31_0_sva_8;
  reg state_3_3_31_0_sva_7;
  reg state_3_3_31_0_sva_6;
  reg state_3_3_31_0_sva_5;
  reg state_3_3_31_0_sva_4;
  reg state_3_3_31_0_sva_3;
  reg state_3_3_31_0_sva_2;
  reg state_3_3_31_0_sva_1;
  reg state_3_3_31_0_sva_0;
  reg state_3_3_63_32_sva_31;
  reg state_3_3_63_32_sva_30;
  reg state_3_3_63_32_sva_29;
  reg state_3_3_63_32_sva_28;
  reg state_3_3_63_32_sva_27;
  reg state_3_3_63_32_sva_26;
  reg state_3_3_63_32_sva_25;
  reg state_3_3_63_32_sva_24;
  reg state_3_3_63_32_sva_23;
  reg state_3_3_63_32_sva_22;
  reg state_3_3_63_32_sva_21;
  reg state_3_3_63_32_sva_20;
  reg state_3_3_63_32_sva_19;
  reg state_3_3_63_32_sva_18;
  reg state_3_3_63_32_sva_17;
  reg state_3_3_63_32_sva_16;
  reg state_3_3_63_32_sva_15;
  reg state_3_3_63_32_sva_14;
  reg state_3_3_63_32_sva_13;
  reg state_3_3_63_32_sva_12;
  reg state_3_3_63_32_sva_11;
  reg state_3_3_63_32_sva_10;
  reg state_3_3_63_32_sva_9;
  reg state_3_3_63_32_sva_8;
  reg state_3_3_63_32_sva_7;
  reg state_3_3_63_32_sva_6;
  reg state_3_3_63_32_sva_5;
  reg state_3_3_63_32_sva_4;
  reg state_3_3_63_32_sva_3;
  reg state_3_3_63_32_sva_2;
  reg state_3_3_63_32_sva_1;
  reg state_3_3_63_32_sva_0;
  reg state_4_3_31_0_sva_31;
  reg state_4_3_31_0_sva_30;
  reg state_4_3_31_0_sva_29;
  reg state_4_3_31_0_sva_28;
  reg state_4_3_31_0_sva_27;
  reg state_4_3_31_0_sva_26;
  reg state_4_3_31_0_sva_25;
  reg state_4_3_31_0_sva_24;
  reg state_4_3_31_0_sva_23;
  reg state_4_3_31_0_sva_22;
  reg state_4_3_31_0_sva_21;
  reg state_4_3_31_0_sva_20;
  reg state_4_3_31_0_sva_19;
  reg state_4_3_31_0_sva_18;
  reg state_4_3_31_0_sva_17;
  reg state_4_3_31_0_sva_16;
  reg state_4_3_31_0_sva_15;
  reg state_4_3_31_0_sva_14;
  reg state_4_3_31_0_sva_13;
  reg state_4_3_31_0_sva_12;
  reg state_4_3_31_0_sva_11;
  reg state_4_3_31_0_sva_10;
  reg state_4_3_31_0_sva_9;
  reg state_4_3_31_0_sva_8;
  reg state_4_3_31_0_sva_7;
  reg state_4_3_31_0_sva_6;
  reg state_4_3_31_0_sva_5;
  reg state_4_3_31_0_sva_4;
  reg state_4_3_31_0_sva_3;
  reg state_4_3_31_0_sva_2;
  reg state_4_3_31_0_sva_1;
  reg state_4_3_31_0_sva_0;
  reg state_4_3_63_32_sva_31;
  reg state_4_3_63_32_sva_30;
  reg state_4_3_63_32_sva_29;
  reg state_4_3_63_32_sva_28;
  reg state_4_3_63_32_sva_27;
  reg state_4_3_63_32_sva_26;
  reg state_4_3_63_32_sva_25;
  reg state_4_3_63_32_sva_24;
  reg state_4_3_63_32_sva_23;
  reg state_4_3_63_32_sva_22;
  reg state_4_3_63_32_sva_21;
  reg state_4_3_63_32_sva_20;
  reg state_4_3_63_32_sva_19;
  reg state_4_3_63_32_sva_18;
  reg state_4_3_63_32_sva_17;
  reg state_4_3_63_32_sva_16;
  reg state_4_3_63_32_sva_15;
  reg state_4_3_63_32_sva_14;
  reg state_4_3_63_32_sva_13;
  reg state_4_3_63_32_sva_12;
  reg state_4_3_63_32_sva_11;
  reg state_4_3_63_32_sva_10;
  reg state_4_3_63_32_sva_9;
  reg state_4_3_63_32_sva_8;
  reg state_4_3_63_32_sva_7;
  reg state_4_3_63_32_sva_6;
  reg state_4_3_63_32_sva_5;
  reg state_4_3_63_32_sva_4;
  reg state_4_3_63_32_sva_3;
  reg state_4_3_63_32_sva_2;
  reg state_4_3_63_32_sva_1;
  reg state_4_3_63_32_sva_0;
  wire plaintext_and_1_ssc;
  reg plaintext_63_32_sva_31;
  reg plaintext_63_32_sva_30;
  reg plaintext_63_32_sva_29;
  reg plaintext_63_32_sva_28;
  reg plaintext_63_32_sva_27;
  reg plaintext_63_32_sva_26;
  reg plaintext_63_32_sva_25;
  reg plaintext_63_32_sva_24;
  reg plaintext_63_32_sva_23;
  reg plaintext_63_32_sva_22;
  reg plaintext_63_32_sva_21;
  reg plaintext_63_32_sva_20;
  reg plaintext_63_32_sva_19;
  reg plaintext_63_32_sva_18;
  reg plaintext_63_32_sva_17;
  reg plaintext_63_32_sva_16;
  reg plaintext_63_32_sva_15;
  reg plaintext_63_32_sva_14;
  reg plaintext_63_32_sva_13;
  reg plaintext_63_32_sva_12;
  reg plaintext_63_32_sva_11;
  reg plaintext_63_32_sva_10;
  reg plaintext_63_32_sva_9;
  reg plaintext_63_32_sva_8;
  reg plaintext_63_32_sva_7;
  reg plaintext_63_32_sva_6;
  reg plaintext_63_32_sva_5;
  reg plaintext_63_32_sva_4;
  reg plaintext_63_32_sva_3;
  reg plaintext_63_32_sva_2;
  reg plaintext_63_32_sva_1;
  reg plaintext_63_32_sva_0;
  wire plaintext_and_ssc;
  reg plaintext_31_0_sva_31;
  reg plaintext_31_0_sva_30;
  reg plaintext_31_0_sva_29;
  reg plaintext_31_0_sva_28;
  reg plaintext_31_0_sva_27;
  reg plaintext_31_0_sva_26;
  reg plaintext_31_0_sva_25;
  reg plaintext_31_0_sva_24;
  reg plaintext_31_0_sva_23;
  reg plaintext_31_0_sva_22;
  reg plaintext_31_0_sva_21;
  reg plaintext_31_0_sva_20;
  reg plaintext_31_0_sva_19;
  reg plaintext_31_0_sva_18;
  reg plaintext_31_0_sva_17;
  reg plaintext_31_0_sva_16;
  reg plaintext_31_0_sva_15;
  reg plaintext_31_0_sva_14;
  reg plaintext_31_0_sva_13;
  reg plaintext_31_0_sva_12;
  reg plaintext_31_0_sva_11;
  reg plaintext_31_0_sva_10;
  reg plaintext_31_0_sva_9;
  reg plaintext_31_0_sva_8;
  reg plaintext_31_0_sva_7;
  reg plaintext_31_0_sva_6;
  reg plaintext_31_0_sva_5;
  reg plaintext_31_0_sva_4;
  reg plaintext_31_0_sva_3;
  reg plaintext_31_0_sva_2;
  reg plaintext_31_0_sva_1;
  reg plaintext_31_0_sva_0;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_31;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_27;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_26;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_25;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_24;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_23;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_22;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_21;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_20;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_19;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_18;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_17;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_16;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_15;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_14;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_13;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_12;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_11;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_10;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_9;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_8;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_7;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_6;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_5;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_4;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_3;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_2;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_1;
  wire Encrypt_Top_sbox_and_cse_63_32_sva_1_0;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_17;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_9;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_8;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_7;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_6;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_5;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_4;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_3;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_2;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_1;
  wire Encrypt_Top_sbox_and_cse_31_0_sva_1_0;
  wire or_2210_cse;
  wire or_1265_cse;
  wire state_and_320_cse;
  wire z_out_1_2;

  wire PLEN_xor_62_nl;
  wire xor_403_nl;
  wire xor_262_nl;
  wire PLEN_xor_60_nl;
  wire xor_418_nl;
  wire xor_260_nl;
  wire PLEN_xor_58_nl;
  wire xor_432_nl;
  wire xor_258_nl;
  wire xor_321_nl;
  wire PLEN_xor_56_nl;
  wire xor_447_nl;
  wire xor_256_nl;
  wire xor_319_nl;
  wire PLEN_xor_54_nl;
  wire xor_462_nl;
  wire xor_254_nl;
  wire xor_317_nl;
  wire PLEN_xor_52_nl;
  wire xor_477_nl;
  wire xor_252_nl;
  wire xor_315_nl;
  wire PLEN_xor_50_nl;
  wire xor_492_nl;
  wire xor_250_nl;
  wire xor_313_nl;
  wire PLEN_xor_48_nl;
  wire xor_506_nl;
  wire xor_248_nl;
  wire xor_311_nl;
  wire PLEN_xor_46_nl;
  wire xor_520_nl;
  wire xor_246_nl;
  wire PLEN_xor_44_nl;
  wire xor_533_nl;
  wire xor_244_nl;
  wire PLEN_xor_42_nl;
  wire xor_546_nl;
  wire xor_242_nl;
  wire xor_305_nl;
  wire PLEN_xor_40_nl;
  wire xor_558_nl;
  wire xor_240_nl;
  wire xor_303_nl;
  wire PLEN_xor_38_nl;
  wire xor_568_nl;
  wire xor_238_nl;
  wire xor_301_nl;
  wire PLEN_xor_36_nl;
  wire xor_579_nl;
  wire xor_236_nl;
  wire xor_299_nl;
  wire PLEN_xor_34_nl;
  wire xor_591_nl;
  wire xor_234_nl;
  wire xor_297_nl;
  wire PLEN_xor_nl;
  wire xor_604_nl;
  wire xor_232_nl;
  wire xor_295_nl;
  wire PLEN_xor_33_nl;
  wire xor_615_nl;
  wire xor_230_nl;
  wire xor_293_nl;
  wire PLEN_xor_35_nl;
  wire xor_626_nl;
  wire xor_228_nl;
  wire xor_291_nl;
  wire PLEN_xor_37_nl;
  wire xor_637_nl;
  wire xor_226_nl;
  wire xor_289_nl;
  wire PLEN_xor_39_nl;
  wire xor_649_nl;
  wire xor_224_nl;
  wire xor_287_nl;
  wire PLEN_xor_41_nl;
  wire xor_660_nl;
  wire xor_222_nl;
  wire xor_285_nl;
  wire PLEN_xor_43_nl;
  wire xor_672_nl;
  wire xor_220_nl;
  wire xor_283_nl;
  wire PLEN_xor_45_nl;
  wire xor_683_nl;
  wire xor_218_nl;
  wire xor_281_nl;
  wire PLEN_xor_47_nl;
  wire xor_692_nl;
  wire xor_216_nl;
  wire xor_279_nl;
  wire PLEN_xor_49_nl;
  wire xor_701_nl;
  wire xor_214_nl;
  wire xor_277_nl;
  wire PLEN_xor_51_nl;
  wire xor_711_nl;
  wire xor_212_nl;
  wire xor_275_nl;
  wire PLEN_xor_53_nl;
  wire xor_721_nl;
  wire xor_210_nl;
  wire xor_316_nl;
  wire xor_273_nl;
  wire PLEN_xor_55_nl;
  wire xor_731_nl;
  wire xor_208_nl;
  wire xor_318_nl;
  wire xor_271_nl;
  wire PLEN_xor_57_nl;
  wire xor_741_nl;
  wire xor_206_nl;
  wire xor_320_nl;
  wire xor_269_nl;
  wire PLEN_xor_59_nl;
  wire xor_751_nl;
  wire xor_204_nl;
  wire xor_322_nl;
  wire xor_267_nl;
  wire PLEN_xor_61_nl;
  wire xor_760_nl;
  wire xor_202_nl;
  wire xor_324_nl;
  wire xor_265_nl;
  wire PLEN_xor_63_nl;
  wire xor_769_nl;
  wire xor_9_nl;
  wire xor_326_nl;
  wire xor_11_nl;
  wire state_xor_338_nl;
  wire state_xor_340_nl;
  wire state_xor_342_nl;
  wire state_xor_344_nl;
  wire state_xor_346_nl;
  wire state_xor_348_nl;
  wire state_xor_350_nl;
  wire state_xor_352_nl;
  wire state_xor_354_nl;
  wire state_xor_356_nl;
  wire state_xor_358_nl;
  wire state_xor_360_nl;
  wire state_xor_362_nl;
  wire state_xor_364_nl;
  wire state_xor_366_nl;
  wire state_xor_368_nl;
  wire state_xor_370_nl;
  wire state_xor_372_nl;
  wire state_xor_374_nl;
  wire state_xor_376_nl;
  wire state_xor_378_nl;
  wire state_xor_380_nl;
  wire state_xor_382_nl;
  wire state_xor_384_nl;
  wire state_xor_386_nl;
  wire state_xor_388_nl;
  wire state_xor_390_nl;
  wire state_xor_392_nl;
  wire state_xor_394_nl;
  wire state_xor_396_nl;
  wire state_xor_398_nl;
  wire state_xor_400_nl;
  wire state_xor_402_nl;
  wire state_xor_404_nl;
  wire state_xor_406_nl;
  wire state_xor_408_nl;
  wire state_xor_410_nl;
  wire state_xor_412_nl;
  wire state_xor_414_nl;
  wire state_xor_416_nl;
  wire state_xor_418_nl;
  wire state_xor_420_nl;
  wire state_xor_422_nl;
  wire state_xor_424_nl;
  wire state_xor_426_nl;
  wire state_xor_428_nl;
  wire state_xor_430_nl;
  wire state_xor_432_nl;
  wire state_xor_434_nl;
  wire state_xor_436_nl;
  wire state_xor_438_nl;
  wire state_xor_440_nl;
  wire state_xor_442_nl;
  wire state_xor_444_nl;
  wire state_xor_446_nl;
  wire state_xor_448_nl;
  wire state_xor_450_nl;
  wire state_xor_452_nl;
  wire state_xor_454_nl;
  wire state_xor_456_nl;
  wire state_xor_458_nl;
  wire state_xor_460_nl;
  wire state_xor_462_nl;
  wire state_xor_464_nl;
  wire state_xor_401_nl;
  wire state_xor_399_nl;
  wire state_xor_397_nl;
  wire state_xor_395_nl;
  wire state_xor_393_nl;
  wire state_xor_391_nl;
  wire state_xor_389_nl;
  wire state_xor_387_nl;
  wire state_xor_385_nl;
  wire state_xor_383_nl;
  wire state_xor_381_nl;
  wire state_xor_379_nl;
  wire state_xor_377_nl;
  wire state_xor_375_nl;
  wire state_xor_373_nl;
  wire state_xor_371_nl;
  wire state_xor_369_nl;
  wire state_xor_367_nl;
  wire state_xor_365_nl;
  wire state_xor_363_nl;
  wire state_xor_361_nl;
  wire state_xor_359_nl;
  wire state_xor_357_nl;
  wire state_xor_355_nl;
  wire state_xor_353_nl;
  wire state_xor_351_nl;
  wire state_xor_349_nl;
  wire state_xor_347_nl;
  wire state_xor_345_nl;
  wire state_xor_343_nl;
  wire state_xor_341_nl;
  wire state_xor_339_nl;
  wire state_xor_465_nl;
  wire state_xor_463_nl;
  wire state_xor_461_nl;
  wire state_xor_459_nl;
  wire state_xor_457_nl;
  wire state_xor_455_nl;
  wire state_xor_453_nl;
  wire state_xor_451_nl;
  wire state_xor_449_nl;
  wire state_xor_447_nl;
  wire state_xor_445_nl;
  wire state_xor_443_nl;
  wire state_xor_441_nl;
  wire state_xor_439_nl;
  wire state_xor_437_nl;
  wire state_xor_435_nl;
  wire state_xor_433_nl;
  wire state_xor_431_nl;
  wire state_xor_429_nl;
  wire state_xor_427_nl;
  wire state_xor_425_nl;
  wire state_xor_423_nl;
  wire state_xor_421_nl;
  wire state_xor_419_nl;
  wire state_xor_417_nl;
  wire state_xor_415_nl;
  wire state_xor_413_nl;
  wire state_xor_411_nl;
  wire state_xor_409_nl;
  wire state_xor_407_nl;
  wire state_xor_405_nl;
  wire state_xor_403_nl;
  wire mux1h_nl;
  wire state_xor_nl;
  wire state_xor_1_nl;
  wire state_xor_2_nl;
  wire state_xor_3_nl;
  wire mux1h_1_nl;
  wire state_xor_4_nl;
  wire state_xor_5_nl;
  wire state_xor_6_nl;
  wire state_xor_7_nl;
  wire mux1h_2_nl;
  wire state_xor_8_nl;
  wire state_xor_9_nl;
  wire state_xor_10_nl;
  wire state_xor_11_nl;
  wire mux1h_3_nl;
  wire state_xor_12_nl;
  wire state_xor_13_nl;
  wire state_xor_14_nl;
  wire state_xor_15_nl;
  wire mux1h_4_nl;
  wire state_xor_16_nl;
  wire state_xor_17_nl;
  wire state_xor_19_nl;
  wire mux1h_5_nl;
  wire state_xor_20_nl;
  wire state_xor_21_nl;
  wire state_xor_23_nl;
  wire mux1h_6_nl;
  wire state_xor_24_nl;
  wire state_xor_25_nl;
  wire state_xor_27_nl;
  wire mux1h_7_nl;
  wire state_xor_28_nl;
  wire state_xor_29_nl;
  wire state_xor_31_nl;
  wire state_xnor_nl;
  wire state_xnor_1_nl;
  wire xor_53_nl;
  wire state_xnor_2_nl;
  wire state_xnor_3_nl;
  wire xor_51_nl;
  wire state_xnor_4_nl;
  wire state_xnor_5_nl;
  wire xor_49_nl;
  wire state_xnor_6_nl;
  wire state_xnor_7_nl;
  wire xor_47_nl;
  wire state_xnor_8_nl;
  wire state_xnor_9_nl;
  wire xor_45_nl;
  wire state_xnor_10_nl;
  wire state_xnor_11_nl;
  wire xor_43_nl;
  wire state_xnor_12_nl;
  wire state_xnor_13_nl;
  wire xor_41_nl;
  wire state_xnor_14_nl;
  wire state_xnor_15_nl;
  wire xor_39_nl;
  wire state_xnor_16_nl;
  wire state_xnor_17_nl;
  wire xor_37_nl;
  wire state_xnor_18_nl;
  wire state_xnor_19_nl;
  wire xor_35_nl;
  wire state_xnor_20_nl;
  wire state_xnor_21_nl;
  wire xor_33_nl;
  wire state_xnor_22_nl;
  wire state_xnor_23_nl;
  wire xor_31_nl;
  wire state_xnor_24_nl;
  wire state_xnor_25_nl;
  wire xor_29_nl;
  wire state_xnor_26_nl;
  wire state_xnor_27_nl;
  wire xor_27_nl;
  wire state_xnor_28_nl;
  wire state_xnor_29_nl;
  wire xor_25_nl;
  wire state_xnor_30_nl;
  wire state_xnor_31_nl;
  wire xor_23_nl;
  wire state_xnor_32_nl;
  wire state_xnor_33_nl;
  wire xor_21_nl;
  wire state_xnor_34_nl;
  wire state_xnor_35_nl;
  wire state_xnor_36_nl;
  wire xor_19_nl;
  wire state_xnor_37_nl;
  wire state_xnor_38_nl;
  wire state_xnor_39_nl;
  wire xor_17_nl;
  wire state_xnor_40_nl;
  wire state_xnor_41_nl;
  wire state_xnor_42_nl;
  wire xor_15_nl;
  wire state_xnor_43_nl;
  wire state_xnor_44_nl;
  wire state_xnor_45_nl;
  wire xor_13_nl;
  wire state_xnor_46_nl;
  wire state_xnor_47_nl;
  wire state_xnor_48_nl;
  wire xor_7_nl;
  wire state_xnor_49_nl;
  wire state_xnor_50_nl;
  wire state_xnor_51_nl;
  wire state_xnor_52_nl;
  wire state_xnor_53_nl;
  wire state_xnor_54_nl;
  wire state_xnor_55_nl;
  wire state_xnor_56_nl;
  wire state_xnor_57_nl;
  wire state_xnor_58_nl;
  wire state_xnor_59_nl;
  wire state_xnor_60_nl;
  wire state_xnor_61_nl;
  wire state_xnor_62_nl;
  wire state_xnor_63_nl;
  wire state_xnor_64_nl;
  wire state_xnor_65_nl;
  wire state_xnor_66_nl;
  wire state_xnor_67_nl;
  wire state_xnor_68_nl;
  wire state_xnor_69_nl;
  wire state_xnor_70_nl;
  wire state_xnor_71_nl;
  wire state_xnor_72_nl;
  wire state_xnor_73_nl;
  wire state_xnor_74_nl;
  wire state_xnor_75_nl;
  wire state_xnor_76_nl;
  wire state_xnor_77_nl;
  wire state_xnor_78_nl;
  wire state_xnor_79_nl;
  wire state_xnor_80_nl;
  wire state_xnor_81_nl;
  wire state_xnor_82_nl;
  wire state_xnor_83_nl;
  wire state_xnor_84_nl;
  wire state_xnor_85_nl;
  wire state_xnor_86_nl;
  wire state_xnor_87_nl;
  wire state_xnor_88_nl;
  wire state_xnor_89_nl;
  wire state_xnor_90_nl;
  wire state_xnor_91_nl;
  wire state_xnor_92_nl;
  wire state_xnor_93_nl;
  wire state_xnor_94_nl;
  wire state_xnor_95_nl;
  wire state_xnor_96_nl;
  wire state_xnor_97_nl;
  wire state_xnor_98_nl;
  wire state_xnor_99_nl;
  wire state_xnor_100_nl;
  wire state_xnor_101_nl;
  wire state_xnor_102_nl;
  wire state_xnor_103_nl;
  wire state_xnor_104_nl;
  wire state_xnor_105_nl;
  wire state_xnor_106_nl;
  wire state_xnor_107_nl;
  wire state_xnor_108_nl;
  wire state_xnor_109_nl;
  wire state_xnor_110_nl;
  wire state_xnor_111_nl;
  wire state_xnor_112_nl;
  wire state_xnor_113_nl;
  wire state_xnor_114_nl;
  wire state_xnor_115_nl;
  wire state_xnor_116_nl;
  wire state_xnor_117_nl;
  wire state_xnor_118_nl;
  wire state_xnor_119_nl;
  wire state_xnor_120_nl;
  wire state_xnor_121_nl;
  wire state_xnor_122_nl;
  wire state_xnor_123_nl;
  wire state_xnor_124_nl;
  wire state_xnor_125_nl;
  wire state_xnor_126_nl;
  wire state_xnor_127_nl;
  wire state_xnor_128_nl;
  wire state_xnor_129_nl;
  wire Encrypt_Top_linear_2_xnor_nl;
  wire xor_64_nl;
  wire state_xnor_130_nl;
  wire state_xnor_131_nl;
  wire state_xnor_132_nl;
  wire Encrypt_Top_linear_2_xnor_1_nl;
  wire xor_66_nl;
  wire state_xnor_133_nl;
  wire state_xnor_134_nl;
  wire state_xnor_135_nl;
  wire Encrypt_Top_linear_2_xnor_2_nl;
  wire xor_68_nl;
  wire state_xnor_136_nl;
  wire state_xnor_137_nl;
  wire state_xnor_138_nl;
  wire Encrypt_Top_linear_2_xnor_3_nl;
  wire xor_70_nl;
  wire state_xnor_139_nl;
  wire state_xnor_140_nl;
  wire state_xnor_141_nl;
  wire Encrypt_Top_linear_2_xnor_4_nl;
  wire xor_72_nl;
  wire state_xnor_142_nl;
  wire state_xnor_143_nl;
  wire state_xnor_144_nl;
  wire Encrypt_Top_linear_2_xnor_5_nl;
  wire xor_74_nl;
  wire state_xnor_145_nl;
  wire state_xnor_146_nl;
  wire state_xnor_147_nl;
  wire state_xnor_148_nl;
  wire state_xnor_149_nl;
  wire state_xnor_150_nl;
  wire state_xnor_151_nl;
  wire mux1h_64_nl;
  wire state_xor_82_nl;
  wire state_xor_83_nl;
  wire state_xor_84_nl;
  wire mux1h_65_nl;
  wire state_xor_85_nl;
  wire state_xor_86_nl;
  wire state_xor_87_nl;
  wire mux1h_66_nl;
  wire state_xor_88_nl;
  wire state_xor_89_nl;
  wire state_xor_90_nl;
  wire mux1h_67_nl;
  wire state_xor_91_nl;
  wire state_xor_92_nl;
  wire state_xor_93_nl;
  wire mux1h_68_nl;
  wire state_xor_94_nl;
  wire state_xor_95_nl;
  wire state_xor_96_nl;
  wire mux1h_69_nl;
  wire state_xor_97_nl;
  wire state_xor_98_nl;
  wire state_xor_99_nl;
  wire mux1h_70_nl;
  wire state_xor_100_nl;
  wire state_xor_101_nl;
  wire state_xor_102_nl;
  wire mux1h_71_nl;
  wire state_xor_103_nl;
  wire state_xor_104_nl;
  wire state_xor_105_nl;
  wire mux1h_72_nl;
  wire state_xor_106_nl;
  wire state_xor_107_nl;
  wire state_xor_108_nl;
  wire mux1h_73_nl;
  wire state_xor_109_nl;
  wire state_xor_110_nl;
  wire state_xor_111_nl;
  wire mux1h_74_nl;
  wire state_xor_112_nl;
  wire state_xor_113_nl;
  wire state_xor_114_nl;
  wire mux1h_75_nl;
  wire state_xor_115_nl;
  wire state_xor_116_nl;
  wire state_xor_117_nl;
  wire mux1h_76_nl;
  wire state_xor_118_nl;
  wire state_xor_119_nl;
  wire state_xor_120_nl;
  wire mux1h_77_nl;
  wire state_xor_121_nl;
  wire state_xor_122_nl;
  wire state_xor_123_nl;
  wire mux1h_78_nl;
  wire state_xor_124_nl;
  wire state_xor_125_nl;
  wire state_xor_126_nl;
  wire mux1h_79_nl;
  wire state_xor_127_nl;
  wire state_xor_128_nl;
  wire state_xor_129_nl;
  wire mux1h_80_nl;
  wire state_xor_130_nl;
  wire state_xor_131_nl;
  wire state_xor_132_nl;
  wire mux1h_81_nl;
  wire state_xor_133_nl;
  wire state_xor_134_nl;
  wire state_xor_135_nl;
  wire mux1h_82_nl;
  wire state_xor_136_nl;
  wire state_xor_137_nl;
  wire state_xor_138_nl;
  wire mux1h_83_nl;
  wire state_xor_139_nl;
  wire state_xor_140_nl;
  wire state_xor_141_nl;
  wire mux1h_84_nl;
  wire state_xor_142_nl;
  wire state_xor_143_nl;
  wire state_xor_144_nl;
  wire mux1h_85_nl;
  wire state_xor_145_nl;
  wire state_xor_146_nl;
  wire state_xor_147_nl;
  wire mux1h_86_nl;
  wire state_xor_148_nl;
  wire state_xor_149_nl;
  wire state_xor_150_nl;
  wire mux1h_87_nl;
  wire state_xor_151_nl;
  wire state_xor_152_nl;
  wire state_xor_153_nl;
  wire mux1h_88_nl;
  wire state_xor_154_nl;
  wire state_xor_155_nl;
  wire state_xor_156_nl;
  wire mux1h_89_nl;
  wire state_xor_157_nl;
  wire state_xor_158_nl;
  wire state_xor_159_nl;
  wire mux1h_90_nl;
  wire state_xor_160_nl;
  wire state_xor_161_nl;
  wire state_xor_162_nl;
  wire state_xor_164_nl;
  wire mux1h_91_nl;
  wire state_xor_165_nl;
  wire state_xor_166_nl;
  wire state_xor_167_nl;
  wire state_xor_169_nl;
  wire mux1h_92_nl;
  wire state_xor_170_nl;
  wire state_xor_171_nl;
  wire state_xor_172_nl;
  wire state_xor_173_nl;
  wire mux1h_93_nl;
  wire state_xor_174_nl;
  wire state_xor_175_nl;
  wire state_xor_176_nl;
  wire state_xor_177_nl;
  wire mux1h_94_nl;
  wire state_xor_178_nl;
  wire state_xor_179_nl;
  wire state_xor_180_nl;
  wire state_xor_181_nl;
  wire mux1h_95_nl;
  wire state_xor_182_nl;
  wire state_xor_183_nl;
  wire state_xor_184_nl;
  wire state_xor_185_nl;
  wire mux1h_96_nl;
  wire state_xor_186_nl;
  wire state_xor_187_nl;
  wire state_xor_188_nl;
  wire state_xor_189_nl;
  wire mux1h_97_nl;
  wire state_xor_190_nl;
  wire state_xor_191_nl;
  wire state_xor_192_nl;
  wire state_xor_193_nl;
  wire mux1h_98_nl;
  wire state_xor_194_nl;
  wire state_xor_195_nl;
  wire state_xor_196_nl;
  wire mux1h_99_nl;
  wire state_xor_197_nl;
  wire state_xor_198_nl;
  wire state_xor_199_nl;
  wire state_xor_200_nl;
  wire mux1h_100_nl;
  wire state_xor_201_nl;
  wire state_xor_202_nl;
  wire state_xor_203_nl;
  wire state_xor_204_nl;
  wire mux1h_101_nl;
  wire state_xor_205_nl;
  wire state_xor_206_nl;
  wire state_xor_207_nl;
  wire state_xor_208_nl;
  wire mux1h_102_nl;
  wire state_xor_209_nl;
  wire state_xor_210_nl;
  wire state_xor_211_nl;
  wire state_xor_212_nl;
  wire mux1h_103_nl;
  wire state_xor_213_nl;
  wire state_xor_214_nl;
  wire state_xor_215_nl;
  wire state_xor_216_nl;
  wire mux1h_104_nl;
  wire state_xor_217_nl;
  wire state_xor_218_nl;
  wire state_xor_219_nl;
  wire state_xor_220_nl;
  wire mux1h_105_nl;
  wire state_xor_221_nl;
  wire state_xor_222_nl;
  wire state_xor_223_nl;
  wire state_xor_224_nl;
  wire mux1h_106_nl;
  wire state_xor_225_nl;
  wire state_xor_226_nl;
  wire state_xor_227_nl;
  wire state_xor_228_nl;
  wire mux1h_107_nl;
  wire state_xor_229_nl;
  wire state_xor_230_nl;
  wire state_xor_231_nl;
  wire mux1h_108_nl;
  wire state_xor_232_nl;
  wire state_xor_233_nl;
  wire state_xor_234_nl;
  wire mux1h_109_nl;
  wire state_xor_235_nl;
  wire state_xor_236_nl;
  wire state_xor_237_nl;
  wire mux1h_110_nl;
  wire state_xor_238_nl;
  wire state_xor_239_nl;
  wire state_xor_240_nl;
  wire mux1h_111_nl;
  wire state_xor_241_nl;
  wire state_xor_242_nl;
  wire state_xor_243_nl;
  wire mux1h_112_nl;
  wire state_xor_244_nl;
  wire state_xor_245_nl;
  wire state_xor_246_nl;
  wire mux1h_113_nl;
  wire state_xor_247_nl;
  wire state_xor_248_nl;
  wire state_xor_249_nl;
  wire mux1h_114_nl;
  wire state_xor_250_nl;
  wire state_xor_251_nl;
  wire state_xor_252_nl;
  wire mux1h_115_nl;
  wire state_xor_253_nl;
  wire state_xor_254_nl;
  wire state_xor_255_nl;
  wire mux1h_116_nl;
  wire state_xor_256_nl;
  wire state_xor_257_nl;
  wire state_xor_258_nl;
  wire mux1h_117_nl;
  wire state_xor_259_nl;
  wire state_xor_260_nl;
  wire state_xor_261_nl;
  wire mux1h_118_nl;
  wire state_xor_262_nl;
  wire state_xor_263_nl;
  wire mux1h_119_nl;
  wire state_xor_264_nl;
  wire state_xor_265_nl;
  wire state_xnor_152_nl;
  wire state_xnor_153_nl;
  wire state_xnor_155_nl;
  wire state_xnor_156_nl;
  wire state_xnor_158_nl;
  wire xor_69_nl;
  wire state_xnor_159_nl;
  wire state_xnor_161_nl;
  wire xor_67_nl;
  wire state_xnor_162_nl;
  wire state_xnor_164_nl;
  wire xor_65_nl;
  wire state_xnor_165_nl;
  wire state_xnor_167_nl;
  wire xor_63_nl;
  wire state_xnor_168_nl;
  wire state_xnor_170_nl;
  wire xor_61_nl;
  wire state_xnor_171_nl;
  wire state_xnor_173_nl;
  wire xor_59_nl;
  wire state_xnor_174_nl;
  wire[3:0] ADLEN_i_ADLEN_i_mux_nl;
  wire nor_28_nl;
  wire state_xor_466_nl;
  wire state_xor_467_nl;
  wire xor_136_nl;
  wire state_xor_468_nl;
  wire state_xor_470_nl;
  wire state_xor_471_nl;
  wire xor_134_nl;
  wire state_xor_472_nl;
  wire state_xor_474_nl;
  wire state_xor_475_nl;
  wire xor_132_nl;
  wire state_xor_476_nl;
  wire state_xor_478_nl;
  wire state_xor_479_nl;
  wire xor_130_nl;
  wire state_xor_480_nl;
  wire state_xor_482_nl;
  wire state_xor_483_nl;
  wire xor_128_nl;
  wire state_xor_484_nl;
  wire state_xor_486_nl;
  wire state_xor_487_nl;
  wire xor_126_nl;
  wire state_xor_488_nl;
  wire state_xor_490_nl;
  wire state_xor_491_nl;
  wire xor_124_nl;
  wire state_xor_492_nl;
  wire state_xor_494_nl;
  wire state_xor_495_nl;
  wire xor_122_nl;
  wire state_xor_496_nl;
  wire state_xor_498_nl;
  wire state_xor_499_nl;
  wire xor_116_nl;
  wire state_xor_500_nl;
  wire state_xor_502_nl;
  wire xor_114_nl;
  wire state_xor_503_nl;
  wire state_xor_505_nl;
  wire xor_112_nl;
  wire state_xor_506_nl;
  wire state_xor_508_nl;
  wire xor_110_nl;
  wire state_xor_509_nl;
  wire state_xor_511_nl;
  wire xor_108_nl;
  wire state_xor_512_nl;
  wire state_xor_514_nl;
  wire xor_106_nl;
  wire state_xor_515_nl;
  wire state_xor_517_nl;
  wire xor_104_nl;
  wire state_xor_518_nl;
  wire state_xor_520_nl;
  wire xor_102_nl;
  wire state_xor_521_nl;
  wire state_xor_523_nl;
  wire xor_100_nl;
  wire state_xor_524_nl;
  wire state_xor_526_nl;
  wire xor_98_nl;
  wire state_xor_527_nl;
  wire state_xor_529_nl;
  wire xor_96_nl;
  wire state_xor_530_nl;
  wire state_xor_532_nl;
  wire xor_94_nl;
  wire state_xor_533_nl;
  wire state_xor_535_nl;
  wire xor_92_nl;
  wire state_xor_536_nl;
  wire state_xor_538_nl;
  wire xor_90_nl;
  wire state_xor_539_nl;
  wire state_xor_541_nl;
  wire xor_88_nl;
  wire state_xor_542_nl;
  wire state_xor_544_nl;
  wire state_xor_545_nl;
  wire xor_86_nl;
  wire state_xor_546_nl;
  wire state_xor_548_nl;
  wire state_xor_549_nl;
  wire xor_84_nl;
  wire state_xor_550_nl;
  wire state_xor_552_nl;
  wire state_xor_553_nl;
  wire xor_82_nl;
  wire state_xor_554_nl;
  wire state_xor_556_nl;
  wire state_xor_557_nl;
  wire xor_80_nl;
  wire state_xor_558_nl;
  wire state_xor_560_nl;
  wire state_xor_561_nl;
  wire xor_78_nl;
  wire state_xor_562_nl;
  wire state_xor_564_nl;
  wire state_xor_565_nl;
  wire xor_76_nl;
  wire state_xor_566_nl;
  wire state_xor_568_nl;
  wire state_xor_569_nl;
  wire xor_5_nl;
  wire state_xor_570_nl;
  wire state_xor_572_nl;
  wire state_xor_573_nl;
  wire xor_75_nl;
  wire state_xor_574_nl;
  wire state_xor_575_nl;
  wire state_xor_576_nl;
  wire xor_77_nl;
  wire state_xor_577_nl;
  wire state_xor_578_nl;
  wire state_xor_579_nl;
  wire xor_79_nl;
  wire state_xor_580_nl;
  wire state_xor_581_nl;
  wire xor_81_nl;
  wire state_xor_582_nl;
  wire state_xor_583_nl;
  wire xor_83_nl;
  wire state_xor_584_nl;
  wire state_xor_585_nl;
  wire xor_85_nl;
  wire state_xor_586_nl;
  wire state_xor_587_nl;
  wire xor_87_nl;
  wire state_xor_588_nl;
  wire state_xor_589_nl;
  wire xor_89_nl;
  wire state_xor_590_nl;
  wire state_xor_591_nl;
  wire xor_91_nl;
  wire state_xor_592_nl;
  wire state_xor_593_nl;
  wire xor_93_nl;
  wire state_xor_594_nl;
  wire state_xor_595_nl;
  wire xor_95_nl;
  wire state_xor_596_nl;
  wire state_xor_597_nl;
  wire xor_97_nl;
  wire state_xor_598_nl;
  wire state_xor_599_nl;
  wire xor_99_nl;
  wire state_xor_600_nl;
  wire state_xor_601_nl;
  wire xor_101_nl;
  wire state_xor_602_nl;
  wire state_xor_603_nl;
  wire xor_103_nl;
  wire state_xor_604_nl;
  wire state_xor_605_nl;
  wire xor_105_nl;
  wire state_xor_606_nl;
  wire state_xor_607_nl;
  wire xor_107_nl;
  wire state_xor_608_nl;
  wire state_xor_609_nl;
  wire xor_109_nl;
  wire state_xor_610_nl;
  wire state_xor_611_nl;
  wire xor_111_nl;
  wire state_xor_612_nl;
  wire state_xor_613_nl;
  wire xor_113_nl;
  wire state_xor_614_nl;
  wire state_xor_615_nl;
  wire xor_115_nl;
  wire state_xor_616_nl;
  wire state_xor_617_nl;
  wire xor_117_nl;
  wire state_xor_618_nl;
  wire state_xor_619_nl;
  wire xor_119_nl;
  wire state_xor_620_nl;
  wire state_xor_621_nl;
  wire xor_121_nl;
  wire state_xor_622_nl;
  wire state_xor_623_nl;
  wire xor_123_nl;
  wire state_xor_624_nl;
  wire state_xor_625_nl;
  wire xor_125_nl;
  wire state_xor_626_nl;
  wire state_xor_627_nl;
  wire xor_127_nl;
  wire state_xor_628_nl;
  wire state_xor_629_nl;
  wire xor_129_nl;
  wire state_xor_630_nl;
  wire state_xor_631_nl;
  wire xor_131_nl;
  wire state_xor_632_nl;
  wire state_xor_633_nl;
  wire xor_133_nl;
  wire state_xor_634_nl;
  wire state_xor_635_nl;
  wire xor_135_nl;
  wire state_xor_636_nl;
  wire state_xor_637_nl;
  wire xor_137_nl;
  wire state_xor_638_nl;
  wire state_xor_639_nl;
  wire xor_120_nl;
  wire state_xor_640_nl;
  wire state_xor_641_nl;
  wire xor_118_nl;
  wire state_xor_642_nl;
  wire state_xor_643_nl;
  wire state_xor_644_nl;
  wire state_xor_645_nl;
  wire state_xor_646_nl;
  wire state_xor_647_nl;
  wire state_xor_648_nl;
  wire state_xor_649_nl;
  wire state_xor_650_nl;
  wire state_xor_651_nl;
  wire state_xor_652_nl;
  wire state_xor_653_nl;
  wire state_xor_654_nl;
  wire state_xor_655_nl;
  wire state_xor_656_nl;
  wire state_xor_657_nl;
  wire state_xor_658_nl;
  wire state_xor_659_nl;
  wire state_xor_660_nl;
  wire state_xor_661_nl;
  wire state_xor_662_nl;
  wire state_xor_663_nl;
  wire state_xor_664_nl;
  wire state_xor_665_nl;
  wire state_xor_666_nl;
  wire state_xor_667_nl;
  wire state_xor_668_nl;
  wire state_xor_670_nl;
  wire state_xor_671_nl;
  wire state_xor_673_nl;
  wire state_xor_674_nl;
  wire state_xor_675_nl;
  wire state_xor_676_nl;
  wire state_xor_677_nl;
  wire state_xor_678_nl;
  wire state_xor_679_nl;
  wire state_xor_680_nl;
  wire state_xor_681_nl;
  wire state_xor_682_nl;
  wire state_xor_683_nl;
  wire state_xor_684_nl;
  wire state_xor_685_nl;
  wire state_xor_686_nl;
  wire state_xor_687_nl;
  wire state_xor_688_nl;
  wire state_xor_689_nl;
  wire state_xor_690_nl;
  wire state_xor_691_nl;
  wire state_xor_692_nl;
  wire state_xor_693_nl;
  wire state_xor_694_nl;
  wire state_xor_695_nl;
  wire state_xor_696_nl;
  wire state_xor_697_nl;
  wire state_xor_698_nl;
  wire state_xor_699_nl;
  wire state_xor_700_nl;
  wire state_xor_701_nl;
  wire state_xor_702_nl;
  wire state_xor_703_nl;
  wire state_xor_704_nl;
  wire state_xor_705_nl;
  wire state_xor_706_nl;
  wire state_xor_707_nl;
  wire state_xor_708_nl;
  wire state_xor_709_nl;
  wire state_xor_710_nl;
  wire state_xor_711_nl;
  wire state_xor_712_nl;
  wire state_xor_713_nl;
  wire state_xor_714_nl;
  wire state_xor_715_nl;
  wire state_xor_716_nl;
  wire state_xor_717_nl;
  wire state_xor_718_nl;
  wire state_xor_719_nl;
  wire state_xor_720_nl;
  wire state_xor_721_nl;
  wire state_xor_722_nl;
  wire state_xor_723_nl;
  wire state_xor_724_nl;
  wire state_xor_725_nl;
  wire state_xor_726_nl;
  wire state_xor_727_nl;
  wire state_xor_728_nl;
  wire state_xor_729_nl;
  wire state_xor_730_nl;
  wire state_xor_731_nl;
  wire state_xor_732_nl;
  wire state_xor_733_nl;
  wire state_xor_734_nl;
  wire state_xor_735_nl;
  wire state_xor_736_nl;
  wire state_xor_737_nl;
  wire state_xor_738_nl;
  wire state_xor_739_nl;
  wire state_xor_740_nl;
  wire state_xor_741_nl;
  wire state_xor_742_nl;
  wire state_xor_743_nl;
  wire state_xor_744_nl;
  wire state_xor_745_nl;
  wire state_xor_746_nl;
  wire state_xor_747_nl;
  wire state_xor_748_nl;
  wire state_xor_749_nl;
  wire state_xor_750_nl;
  wire state_xor_751_nl;
  wire state_xor_752_nl;
  wire state_xor_753_nl;
  wire state_xor_754_nl;
  wire state_xor_755_nl;
  wire state_xor_756_nl;
  wire state_xor_757_nl;
  wire state_xor_758_nl;
  wire state_xor_759_nl;
  wire state_xor_760_nl;
  wire state_xor_761_nl;
  wire state_xor_762_nl;
  wire state_xor_763_nl;
  wire state_xor_764_nl;
  wire state_xor_765_nl;
  wire state_xor_766_nl;
  wire state_xor_767_nl;
  wire state_xor_768_nl;
  wire state_xor_769_nl;
  wire state_xor_770_nl;
  wire state_xor_771_nl;
  wire state_xor_772_nl;
  wire state_xor_773_nl;
  wire state_xor_774_nl;
  wire state_xor_775_nl;
  wire state_xor_776_nl;
  wire state_xor_777_nl;
  wire state_xor_778_nl;
  wire state_xor_779_nl;
  wire state_xor_780_nl;
  wire state_xor_781_nl;
  wire state_xor_782_nl;
  wire state_xor_783_nl;
  wire state_xor_784_nl;
  wire state_xor_785_nl;
  wire state_xor_786_nl;
  wire state_xor_787_nl;
  wire state_xor_788_nl;
  wire state_xor_789_nl;
  wire state_xor_790_nl;
  wire state_xor_791_nl;
  wire state_xor_792_nl;
  wire state_xor_793_nl;
  wire state_xor_794_nl;
  wire state_xor_795_nl;
  wire state_xor_796_nl;
  wire state_xor_797_nl;
  wire state_xor_798_nl;
  wire state_xor_799_nl;
  wire state_xor_800_nl;
  wire state_xor_801_nl;
  wire state_xor_802_nl;
  wire state_xor_803_nl;
  wire state_xor_804_nl;
  wire state_xor_805_nl;
  wire state_xor_806_nl;
  wire state_xor_807_nl;
  wire state_xor_808_nl;
  wire state_xor_809_nl;
  wire state_xor_810_nl;
  wire state_xor_811_nl;
  wire state_xor_812_nl;
  wire state_xor_813_nl;
  wire state_xor_814_nl;
  wire state_xor_815_nl;
  wire state_xor_816_nl;
  wire state_xor_817_nl;
  wire state_xor_818_nl;
  wire state_xor_819_nl;
  wire state_xor_820_nl;
  wire state_xor_821_nl;
  wire state_xor_822_nl;
  wire state_xor_823_nl;
  wire state_xor_824_nl;
  wire state_xor_825_nl;
  wire state_xor_826_nl;
  wire state_xor_827_nl;
  wire state_xor_828_nl;
  wire state_xor_829_nl;
  wire state_xor_830_nl;
  wire state_xor_831_nl;
  wire state_xor_832_nl;
  wire state_xor_833_nl;
  wire state_xor_834_nl;
  wire state_xor_835_nl;
  wire state_xor_836_nl;
  wire state_xor_837_nl;
  wire state_xor_838_nl;
  wire state_xor_839_nl;
  wire state_xor_840_nl;
  wire state_xor_842_nl;
  wire state_xor_843_nl;
  wire state_xor_845_nl;
  wire state_xor_846_nl;
  wire state_xor_848_nl;
  wire state_xor_849_nl;
  wire state_xor_851_nl;
  wire state_xor_852_nl;
  wire state_xor_854_nl;
  wire state_xor_855_nl;
  wire state_xor_857_nl;
  wire state_xor_858_nl;
  wire state_xor_859_nl;
  wire state_xor_860_nl;
  wire state_xor_861_nl;
  wire state_xor_862_nl;
  wire state_xor_863_nl;
  wire state_xor_864_nl;
  wire state_xor_865_nl;
  wire state_xor_866_nl;
  wire state_xor_867_nl;
  wire state_xor_868_nl;
  wire state_xor_869_nl;
  wire state_xor_870_nl;
  wire state_xor_871_nl;
  wire state_xor_872_nl;
  wire state_xor_873_nl;
  wire state_xor_874_nl;
  wire state_xor_875_nl;
  wire state_xor_876_nl;
  wire state_xor_877_nl;
  wire state_xor_878_nl;
  wire state_xor_879_nl;
  wire state_xor_880_nl;
  wire state_xor_881_nl;
  wire state_xor_882_nl;
  wire state_xor_883_nl;
  wire state_xor_884_nl;
  wire state_xor_885_nl;
  wire state_xor_886_nl;
  wire state_xor_887_nl;
  wire state_xor_888_nl;
  wire state_xor_889_nl;
  wire state_xor_890_nl;
  wire state_xor_891_nl;
  wire state_xor_892_nl;
  wire state_xor_893_nl;
  wire state_xor_894_nl;
  wire state_xor_895_nl;
  wire state_xor_896_nl;
  wire state_xor_897_nl;
  wire state_xor_898_nl;
  wire state_xor_899_nl;
  wire state_xor_900_nl;
  wire state_xor_901_nl;
  wire state_xor_902_nl;
  wire state_xor_903_nl;
  wire state_xor_904_nl;
  wire state_xor_905_nl;
  wire state_xor_906_nl;
  wire state_xor_907_nl;
  wire state_xor_908_nl;
  wire state_xor_909_nl;
  wire state_xor_910_nl;
  wire state_xor_911_nl;
  wire state_xor_912_nl;
  wire state_xor_913_nl;
  wire state_xor_914_nl;
  wire state_xor_915_nl;
  wire state_xor_916_nl;
  wire state_xor_917_nl;
  wire state_xor_918_nl;
  wire state_xor_919_nl;
  wire state_xor_920_nl;
  wire state_xor_921_nl;
  wire state_xor_922_nl;
  wire state_xor_923_nl;
  wire state_xor_924_nl;
  wire state_xor_925_nl;
  wire state_xor_926_nl;
  wire state_xor_927_nl;
  wire state_xor_928_nl;
  wire state_xor_929_nl;
  wire state_xor_930_nl;
  wire state_xor_931_nl;
  wire state_xor_932_nl;
  wire state_xor_933_nl;
  wire state_xor_934_nl;
  wire state_xor_935_nl;
  wire state_xor_936_nl;
  wire state_xor_937_nl;
  wire state_xor_938_nl;
  wire state_xor_939_nl;
  wire state_xor_940_nl;
  wire state_xor_941_nl;
  wire state_xor_942_nl;
  wire state_xor_943_nl;
  wire state_xor_944_nl;
  wire state_xor_945_nl;
  wire state_xor_946_nl;
  wire state_xor_947_nl;
  wire state_xor_948_nl;
  wire state_xor_949_nl;
  wire state_xor_950_nl;
  wire state_xor_951_nl;
  wire state_xor_952_nl;
  wire state_xor_953_nl;
  wire state_xor_954_nl;
  wire state_xnor_176_nl;
  wire state_xnor_177_nl;
  wire state_xnor_178_nl;
  wire state_xnor_179_nl;
  wire state_xnor_180_nl;
  wire state_xnor_181_nl;
  wire state_xnor_182_nl;
  wire state_xnor_183_nl;
  wire[7:0] operator_8_false_mux_1_nl;
  wire[2:0] AD_P6_acc_nl;
  wire[3:0] nl_AD_P6_acc_nl;
  wire[1:0] AD_P6_mux_2_nl;
  wire[2:0] INIT_P12_mux_2_nl;
  wire or_2257_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[2:0] AD_P6_acc_4_nl;
  wire[3:0] nl_AD_P6_acc_4_nl;
  wire [3:0] nl_U_ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_rg_I_1;
  assign nl_AD_P6_acc_4_nl = conv_u2u_2_3(AD_P6_j_2_0_sva[2:1]) + 3'b011;
  assign AD_P6_acc_4_nl = nl_AD_P6_acc_4_nl[2:0];
  assign nl_U_ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_rg_I_1 = {AD_P6_acc_4_nl
      , (AD_P6_j_2_0_sva[0])};
  wire [31:0] nl_Encrypt_Top_run_data_out_rsci_inst_data_out_rsci_idat;
  assign nl_Encrypt_Top_run_data_out_rsci_inst_data_out_rsci_idat = {data_out_rsci_idat_31
      , data_out_rsci_idat_30 , data_out_rsci_idat_29 , data_out_rsci_idat_28 , data_out_rsci_idat_27
      , data_out_rsci_idat_26 , data_out_rsci_idat_25 , data_out_rsci_idat_24 , data_out_rsci_idat_23
      , data_out_rsci_idat_22 , data_out_rsci_idat_21 , data_out_rsci_idat_20 , data_out_rsci_idat_19
      , data_out_rsci_idat_18 , data_out_rsci_idat_17 , data_out_rsci_idat_16 , data_out_rsci_idat_15
      , data_out_rsci_idat_14 , data_out_rsci_idat_13 , data_out_rsci_idat_12 , data_out_rsci_idat_11
      , data_out_rsci_idat_10 , data_out_rsci_idat_9 , data_out_rsci_idat_8 , data_out_rsci_idat_7
      , data_out_rsci_idat_6 , data_out_rsci_idat_5 , data_out_rsci_idat_4 , data_out_rsci_idat_3
      , data_out_rsci_idat_2 , data_out_rsci_idat_1 , data_out_rsci_idat_0};
  wire  nl_Encrypt_Top_run_run_fsm_inst_INIT_P12_C_0_tr0;
  assign nl_Encrypt_Top_run_run_fsm_inst_INIT_P12_C_0_tr0 = ~ z_out_1_2;
  wire  nl_Encrypt_Top_run_run_fsm_inst_AD_P6_C_0_tr0;
  assign nl_Encrypt_Top_run_run_fsm_inst_AD_P6_C_0_tr0 = ~ z_out_1_2;
  wire  nl_Encrypt_Top_run_run_fsm_inst_ADLEN_C_2_tr0;
  assign nl_Encrypt_Top_run_run_fsm_inst_ADLEN_C_2_tr0 = (z_out_2[7]) | ((({ADLEN_i_7_0_sva_6_4
      , ADLEN_i_7_0_sva_3_0}) == (z_out[6:0])) & (z_out[8:7]==2'b00));
  wire  nl_Encrypt_Top_run_run_fsm_inst_ENC_P6_C_0_tr0;
  assign nl_Encrypt_Top_run_run_fsm_inst_ENC_P6_C_0_tr0 = ~ z_out_1_2;
  wire  nl_Encrypt_Top_run_run_fsm_inst_FINAL_P12_C_0_tr0;
  assign nl_Encrypt_Top_run_run_fsm_inst_FINAL_P12_C_0_tr0 = ~ z_out_1_2;
  ROM_1i4_1o8_0bc064f669c474330176c941c6dd719bb8  U_ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_rg
      (
      .I_1(ADLEN_i_7_0_sva_3_0),
      .O_1(ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1)
    );
  ROM_1i4_1o8_6f8a8acefa07ca761551b27c9076176eb8  U_ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_rg
      (
      .I_1(nl_U_ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_rg_I_1[3:0]),
      .O_1(ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1)
    );
  Encrypt_Top_run_data_in_rsci Encrypt_Top_run_data_in_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .data_in_rsc_dat(data_in_rsc_dat),
      .data_in_rsc_vld(data_in_rsc_vld),
      .data_in_rsc_rdy(data_in_rsc_rdy),
      .run_wen(run_wen),
      .data_in_rsci_oswt(reg_data_in_rsci_iswt0_cse),
      .data_in_rsci_wen_comp(data_in_rsci_wen_comp),
      .data_in_rsci_idat_mxwt(data_in_rsci_idat_mxwt)
    );
  Encrypt_Top_run_data_out_rsci Encrypt_Top_run_data_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .data_out_rsc_dat(data_out_rsc_dat),
      .data_out_rsc_vld(data_out_rsc_vld),
      .data_out_rsc_rdy(data_out_rsc_rdy),
      .run_wen(run_wen),
      .data_out_rsci_oswt(reg_data_out_rsci_iswt0_cse),
      .data_out_rsci_wen_comp(data_out_rsci_wen_comp),
      .data_out_rsci_idat(nl_Encrypt_Top_run_data_out_rsci_inst_data_out_rsci_idat[31:0])
    );
  Encrypt_Top_run_staller Encrypt_Top_run_staller_inst (
      .run_wen(run_wen),
      .data_in_rsci_wen_comp(data_in_rsci_wen_comp),
      .data_out_rsci_wen_comp(data_out_rsci_wen_comp)
    );
  Encrypt_Top_run_run_fsm Encrypt_Top_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .INIT_P12_C_0_tr0(nl_Encrypt_Top_run_run_fsm_inst_INIT_P12_C_0_tr0),
      .AD_P6_C_0_tr0(nl_Encrypt_Top_run_run_fsm_inst_AD_P6_C_0_tr0),
      .ADLEN_C_2_tr0(nl_Encrypt_Top_run_run_fsm_inst_ADLEN_C_2_tr0),
      .ENC_P6_C_0_tr0(nl_Encrypt_Top_run_run_fsm_inst_ENC_P6_C_0_tr0),
      .PLEN_C_3_tr0(or_dcpl_9),
      .FINAL_P12_C_0_tr0(nl_Encrypt_Top_run_run_fsm_inst_FINAL_P12_C_0_tr0)
    );
  assign or_2210_cse = (fsm_output[7:6]!=2'b00) | and_90_cse | (fsm_output[12]) |
      and_94_cse | (fsm_output[17:15]!=3'b000);
  assign and_4636_cse = run_wen & or_2210_cse;
  assign xor_2168_cse = xor_cse_948 ^ xor_cse_2005;
  assign xor_2162_cse = xor_cse_859 ^ xor_cse_2040;
  assign xor_2172_cse = xor_cse_446 ^ xor_cse_2017;
  assign xor_2184_cse = xor_cse_401 ^ xor_cse_1995;
  assign xor_2186_cse = xor_cse_888 ^ xor_cse_2044;
  assign xor_2182_cse = xor_cse_878 ^ xor_cse_2053;
  assign state_and_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[4]) | (fsm_output[11]) | (fsm_output[13]) | (fsm_output[14]));
  assign state_and_4_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | (fsm_output[4]) | and_21_cse | and_90_cse | (fsm_output[14:13]!=2'b00));
  assign state_and_8_cse = run_wen & ((fsm_output[1:0]!=2'b00) | or_tmp_382 | and_885_cse
      | and_94_cse);
  assign state_and_24_cse = run_wen & ((fsm_output[1:0]!=2'b00) | and_24_cse | and_885_cse
      | and_39_cse | and_94_cse);
  assign state_and_56_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[4])
      | (fsm_output[11]) | and_885_cse | (fsm_output[14]));
  assign state_and_64_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | and_24_cse | (fsm_output[14:13]!=2'b00));
  assign state_and_86_cse = run_wen & ((fsm_output[2:0]!=3'b000) | or_tmp_913 | and_90_cse
      | (fsm_output[14:13]!=2'b00));
  assign state_and_90_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2])
      | (fsm_output[4]) | and_21_cse | and_90_cse | (fsm_output[14:13]!=2'b00));
  assign state_and_92_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[2])
      | (fsm_output[4]) | and_21_cse | and_90_cse | (fsm_output[14]));
  assign state_and_98_cse = run_wen & ((fsm_output[2:0]!=3'b000) | or_tmp_913 | and_90_cse
      | (fsm_output[14]));
  assign state_and_118_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[3])
      | or_tmp_913 | and_90_cse | (fsm_output[14:13]!=2'b00));
  assign state_and_120_cse = run_wen & ((fsm_output[0]) | (fsm_output[1]) | (fsm_output[4])
      | (fsm_output[5]) | (fsm_output[13]) | and_39_cse | and_94_cse);
  assign plaintext_and_ssc = run_wen & ((fsm_output[10]) | (fsm_output[0]) | (fsm_output[1]));
  assign and_21_cse = z_out_1_2 & (fsm_output[11]);
  assign plaintext_and_1_ssc = run_wen & (fsm_output[11:10]==2'b00);
  assign and_39_cse = z_out_1_2 & (fsm_output[14]);
  assign ADLEN_i_and_ssc = run_wen & (and_740_cse | and_738_cse | (fsm_output[5])
      | (fsm_output[8]) | ADLEN_i_7_0_sva_6_0_mx0c3);
  assign or_1265_cse = (fsm_output[14]) | (fsm_output[1]);
  assign state_and_128_cse = run_wen & ((fsm_output[1]) | (fsm_output[4]) | (fsm_output[11])
      | and_885_cse | and_39_cse | and_94_cse);
  assign state_and_137_cse = run_wen & ((fsm_output[1]) | and_24_cse | and_885_cse
      | and_39_cse | and_94_cse);
  assign state_and_158_cse = run_wen & ((fsm_output[1]) | (fsm_output[4]) | (fsm_output[11])
      | and_885_cse | (fsm_output[14]));
  assign state_and_161_cse = run_wen & ((fsm_output[1]) | and_24_cse | and_885_cse
      | (fsm_output[14]));
  assign state_and_192_cse = run_wen & ((fsm_output[1]) | (fsm_output[4]) | (fsm_output[11])
      | (fsm_output[14]));
  assign state_and_201_cse = run_wen & ((fsm_output[1]) | and_24_cse | (fsm_output[14]));
  assign state_and_208_cse = run_wen & ((fsm_output[1]) | or_tmp_1693);
  assign state_and_320_cse = run_wen & ((fsm_output[2]) | (fsm_output[3]) | (fsm_output[18])
      | (fsm_output[17]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]) |
      (fsm_output[11]) | (fsm_output[14]));
  assign ADLEN_ADLEN_xor_2_itm_mx0w0 = (data_in_rsci_idat_mxwt[0]) ^ state_0_32_lpi_6;
  assign state_0_0_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[0]) ^ state_0_0_lpi_6;
  assign data_out_rsci_idat_0_mx0w6 = state_2_32_1_lpi_4 ^ (key3[0]);
  assign data_out_rsci_idat_0_mx0w7 = state_2_0_1_lpi_6 ^ (key4[0]);
  assign ADLEN_ADLEN_xor_4_itm_mx0w0 = (data_in_rsci_idat_mxwt[1]) ^ state_0_33_lpi_6;
  assign state_0_1_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[1]) ^ state_0_1_lpi_6;
  assign data_out_rsci_idat_1_mx0w6 = state_2_33_1_lpi_4 ^ (key3[1]);
  assign data_out_rsci_idat_1_mx0w7 = state_2_1_1_lpi_6 ^ (key4[1]);
  assign ADLEN_ADLEN_xor_6_itm_mx0w0 = (data_in_rsci_idat_mxwt[2]) ^ state_0_34_lpi_6;
  assign state_0_2_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[2]) ^ state_0_2_lpi_6;
  assign data_out_rsci_idat_2_mx0w6 = state_2_34_1_lpi_4 ^ (key3[2]);
  assign ADLEN_ADLEN_xor_8_itm_mx0w0 = (data_in_rsci_idat_mxwt[3]) ^ state_0_35_lpi_6;
  assign state_0_3_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[3]) ^ state_0_3_lpi_6;
  assign data_out_rsci_idat_3_mx0w6 = state_2_35_1_lpi_4 ^ (key3[3]);
  assign ADLEN_ADLEN_xor_10_itm_mx0w0 = (data_in_rsci_idat_mxwt[4]) ^ state_0_36_lpi_6;
  assign state_0_4_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[4]) ^ state_0_4_lpi_6;
  assign data_out_rsci_idat_4_mx0w6 = state_2_36_1_lpi_4 ^ (key3[4]);
  assign ADLEN_ADLEN_xor_12_itm_mx0w0 = (data_in_rsci_idat_mxwt[5]) ^ state_0_37_lpi_6;
  assign state_0_5_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[5]) ^ state_0_5_lpi_6;
  assign data_out_rsci_idat_5_mx0w6 = state_2_37_1_lpi_4 ^ (key3[5]);
  assign ADLEN_ADLEN_xor_14_itm_mx0w0 = (data_in_rsci_idat_mxwt[6]) ^ state_0_38_lpi_6;
  assign state_0_6_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[6]) ^ state_0_6_lpi_6;
  assign data_out_rsci_idat_6_mx0w6 = state_2_38_1_lpi_4 ^ (key3[6]);
  assign ADLEN_ADLEN_xor_16_itm_mx0w0 = (data_in_rsci_idat_mxwt[7]) ^ state_0_39_lpi_6;
  assign state_0_7_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[7]) ^ state_0_7_lpi_6;
  assign data_out_rsci_idat_7_mx0w6 = state_2_39_1_lpi_4 ^ (key3[7]);
  assign ADLEN_ADLEN_xor_18_itm_mx0w0 = (data_in_rsci_idat_mxwt[8]) ^ state_0_40_lpi_6;
  assign state_0_8_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[8]) ^ state_0_8_lpi_6;
  assign data_out_rsci_idat_8_mx0w6 = state_2_40_1_lpi_4 ^ (key3[8]);
  assign data_out_rsci_idat_8_mx0w7 = state_2_8_1_lpi_4 ^ (key4[8]);
  assign ADLEN_ADLEN_xor_20_itm_mx0w0 = (data_in_rsci_idat_mxwt[9]) ^ state_0_41_lpi_6;
  assign state_0_9_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[9]) ^ state_0_9_lpi_6;
  assign data_out_rsci_idat_9_mx0w6 = state_2_41_1_lpi_4 ^ (key3[9]);
  assign data_out_rsci_idat_9_mx0w7 = state_2_9_1_lpi_4 ^ (key4[9]);
  assign ADLEN_ADLEN_xor_22_itm_mx0w0 = (data_in_rsci_idat_mxwt[10]) ^ state_0_42_lpi_6;
  assign state_0_10_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[10]) ^ state_0_10_lpi_6;
  assign data_out_rsci_idat_10_mx0w6 = state_2_42_1_lpi_4 ^ (key3[10]);
  assign ADLEN_ADLEN_xor_24_itm_mx0w0 = (data_in_rsci_idat_mxwt[11]) ^ state_0_43_lpi_6;
  assign state_0_11_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[11]) ^ state_0_11_lpi_6;
  assign data_out_rsci_idat_11_mx0w6 = state_2_43_1_lpi_4 ^ (key3[11]);
  assign ADLEN_ADLEN_xor_26_itm_mx0w0 = (data_in_rsci_idat_mxwt[12]) ^ state_0_44_lpi_6;
  assign state_0_12_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[12]) ^ state_0_12_lpi_6;
  assign data_out_rsci_idat_12_mx0w6 = state_2_44_1_lpi_4 ^ (key3[12]);
  assign ADLEN_ADLEN_xor_28_itm_mx0w0 = (data_in_rsci_idat_mxwt[13]) ^ state_0_45_lpi_6;
  assign state_0_13_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[13]) ^ state_0_13_lpi_6;
  assign data_out_rsci_idat_13_mx0w6 = state_2_45_1_lpi_4 ^ (key3[13]);
  assign ADLEN_ADLEN_xor_30_itm_mx0w0 = (data_in_rsci_idat_mxwt[14]) ^ state_0_46_lpi_6;
  assign state_0_14_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[14]) ^ state_0_14_lpi_6;
  assign data_out_rsci_idat_14_mx0w6 = state_2_46_1_lpi_4 ^ (key3[14]);
  assign ADLEN_ADLEN_xor_32_itm_mx0w0 = (data_in_rsci_idat_mxwt[15]) ^ state_0_47_lpi_6;
  assign state_0_15_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[15]) ^ state_0_15_lpi_6;
  assign data_out_rsci_idat_15_mx0w6 = state_2_47_1_lpi_4 ^ (key3[15]);
  assign ADLEN_ADLEN_xor_34_itm_mx0w0 = (data_in_rsci_idat_mxwt[16]) ^ state_0_48_lpi_6;
  assign state_0_16_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[16]) ^ state_0_16_lpi_6;
  assign data_out_rsci_idat_16_mx0w6 = state_2_48_1_lpi_4 ^ (key3[16]);
  assign ADLEN_ADLEN_xor_36_itm_mx0w0 = (data_in_rsci_idat_mxwt[17]) ^ state_0_49_lpi_6;
  assign state_0_17_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[17]) ^ state_0_17_lpi_6;
  assign data_out_rsci_idat_17_mx0w6 = state_2_49_1_lpi_4 ^ (key3[17]);
  assign ADLEN_ADLEN_xor_38_itm_mx0w0 = (data_in_rsci_idat_mxwt[18]) ^ state_0_50_lpi_6;
  assign state_0_18_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[18]) ^ state_0_18_lpi_6;
  assign data_out_rsci_idat_18_mx0w6 = state_2_50_1_lpi_4 ^ (key3[18]);
  assign ADLEN_ADLEN_xor_40_itm_mx0w0 = (data_in_rsci_idat_mxwt[19]) ^ state_0_51_lpi_6;
  assign state_0_19_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[19]) ^ state_0_19_lpi_6;
  assign data_out_rsci_idat_19_mx0w6 = state_2_51_1_lpi_4 ^ (key3[19]);
  assign ADLEN_ADLEN_xor_42_itm_mx0w0 = (data_in_rsci_idat_mxwt[20]) ^ state_0_52_lpi_6;
  assign state_0_20_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[20]) ^ state_0_20_lpi_6;
  assign data_out_rsci_idat_20_mx0w6 = state_2_52_1_lpi_4 ^ (key3[20]);
  assign ADLEN_ADLEN_xor_44_itm_mx0w0 = (data_in_rsci_idat_mxwt[21]) ^ state_0_53_lpi_6;
  assign state_0_21_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[21]) ^ state_0_21_lpi_6;
  assign data_out_rsci_idat_21_mx0w6 = state_2_53_1_lpi_4 ^ (key3[21]);
  assign ADLEN_ADLEN_xor_46_itm_mx0w0 = (data_in_rsci_idat_mxwt[22]) ^ state_0_54_lpi_6;
  assign state_0_22_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[22]) ^ state_0_22_lpi_6;
  assign data_out_rsci_idat_22_mx0w6 = state_2_54_1_lpi_4 ^ (key3[22]);
  assign ADLEN_ADLEN_xor_48_itm_mx0w0 = (data_in_rsci_idat_mxwt[23]) ^ state_0_55_lpi_6;
  assign state_0_23_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[23]) ^ state_0_23_lpi_6;
  assign data_out_rsci_idat_23_mx0w6 = state_2_55_1_lpi_4 ^ (key3[23]);
  assign ADLEN_ADLEN_xor_50_itm_mx0w0 = (data_in_rsci_idat_mxwt[24]) ^ state_0_56_lpi_6;
  assign state_0_24_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[24]) ^ state_0_24_lpi_6;
  assign data_out_rsci_idat_24_mx0w6 = state_2_56_1_lpi_4 ^ (key3[24]);
  assign ADLEN_ADLEN_xor_52_itm_mx0w0 = (data_in_rsci_idat_mxwt[25]) ^ state_0_57_lpi_6;
  assign state_0_25_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[25]) ^ state_0_25_lpi_6;
  assign data_out_rsci_idat_25_mx0w6 = state_2_57_1_lpi_4 ^ (key3[25]);
  assign ADLEN_ADLEN_xor_54_itm_mx0w0 = (data_in_rsci_idat_mxwt[26]) ^ state_0_58_lpi_6;
  assign state_0_26_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[26]) ^ state_0_26_lpi_6;
  assign ADLEN_ADLEN_xor_56_itm_mx0w0 = (data_in_rsci_idat_mxwt[27]) ^ state_0_59_lpi_6;
  assign state_0_27_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[27]) ^ state_0_27_lpi_6;
  assign ADLEN_ADLEN_xor_58_itm_mx0w0 = (data_in_rsci_idat_mxwt[28]) ^ state_0_60_lpi_6;
  assign state_0_28_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[28]) ^ state_0_28_lpi_6;
  assign ADLEN_ADLEN_xor_60_itm_mx0w0 = (data_in_rsci_idat_mxwt[29]) ^ state_0_61_lpi_6;
  assign state_0_29_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[29]) ^ state_0_29_lpi_6;
  assign ADLEN_ADLEN_xor_62_itm_mx0w0 = (data_in_rsci_idat_mxwt[30]) ^ state_0_62_lpi_6;
  assign state_0_30_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[30]) ^ state_0_30_lpi_6;
  assign ADLEN_ADLEN_xor_64_itm_mx0w0 = (data_in_rsci_idat_mxwt[31]) ^ state_0_63_lpi_6;
  assign state_0_31_sva_2_mx0w1 = (data_in_rsci_idat_mxwt[31]) ^ state_0_31_lpi_6;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_31 = state_4_3_63_32_sva_31 & plaintext_63_32_sva_31;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_27 = state_4_3_63_32_sva_27 & plaintext_63_32_sva_27;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_26 = state_4_3_63_32_sva_26 & plaintext_63_32_sva_26;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_25 = state_4_3_63_32_sva_25 & plaintext_63_32_sva_25;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_24 = state_4_3_63_32_sva_24 & plaintext_63_32_sva_24;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_23 = state_4_3_63_32_sva_23 & plaintext_63_32_sva_23;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_22 = state_4_3_63_32_sva_22 & plaintext_63_32_sva_22;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_21 = state_4_3_63_32_sva_21 & plaintext_63_32_sva_21;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_20 = state_4_3_63_32_sva_20 & plaintext_63_32_sva_20;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_19 = state_4_3_63_32_sva_19 & plaintext_63_32_sva_19;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_18 = state_4_3_63_32_sva_18 & plaintext_63_32_sva_18;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_17 = state_4_3_63_32_sva_17 & plaintext_63_32_sva_17;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_16 = state_4_3_63_32_sva_16 & plaintext_63_32_sva_16;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_15 = state_4_3_63_32_sva_15 & plaintext_63_32_sva_15;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_14 = state_4_3_63_32_sva_14 & plaintext_63_32_sva_14;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_13 = state_4_3_63_32_sva_13 & plaintext_63_32_sva_13;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_12 = state_4_3_63_32_sva_12 & plaintext_63_32_sva_12;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_11 = state_4_3_63_32_sva_11 & plaintext_63_32_sva_11;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_10 = state_4_3_63_32_sva_10 & plaintext_63_32_sva_10;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_9 = state_4_3_63_32_sva_9 & plaintext_63_32_sva_9;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_8 = state_4_3_63_32_sva_8 & plaintext_63_32_sva_8;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_7 = state_4_3_63_32_sva_7 & plaintext_63_32_sva_7;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_6 = state_4_3_63_32_sva_6 & plaintext_63_32_sva_6;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_5 = state_4_3_63_32_sva_5 & plaintext_63_32_sva_5;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_4 = state_4_3_63_32_sva_4 & plaintext_63_32_sva_4;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_3 = state_4_3_63_32_sva_3 & plaintext_63_32_sva_3;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_2 = state_4_3_63_32_sva_2 & plaintext_63_32_sva_2;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_1 = state_4_3_63_32_sva_1 & plaintext_63_32_sva_1;
  assign Encrypt_Top_sbox_and_cse_63_32_sva_1_0 = state_4_3_63_32_sva_0 & plaintext_63_32_sva_0;
  assign Encrypt_Top_sbox_and_2_cse_63_sva_1 = plaintext_63_32_sva_31 & state_0_63_lpi_6;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_17 = state_4_3_31_0_sva_17 & plaintext_31_0_sva_17;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_9 = state_4_3_31_0_sva_9 & plaintext_31_0_sva_9;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_8 = state_4_3_31_0_sva_8 & plaintext_31_0_sva_8;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_7 = state_4_3_31_0_sva_7 & plaintext_31_0_sva_7;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_6 = state_4_3_31_0_sva_6 & plaintext_31_0_sva_6;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_5 = state_4_3_31_0_sva_5 & plaintext_31_0_sva_5;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_4 = state_4_3_31_0_sva_4 & plaintext_31_0_sva_4;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_3 = state_4_3_31_0_sva_3 & plaintext_31_0_sva_3;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_2 = state_4_3_31_0_sva_2 & plaintext_31_0_sva_2;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_1 = state_4_3_31_0_sva_1 & plaintext_31_0_sva_1;
  assign Encrypt_Top_sbox_and_cse_31_0_sva_1_0 = state_4_3_31_0_sva_0 & plaintext_31_0_sva_0;
  assign Encrypt_Top_sbox_and_2_cse_0_sva_1 = plaintext_31_0_sva_0 & state_0_0_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_1_sva_1 = plaintext_31_0_sva_1 & state_0_1_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_2_sva_1 = plaintext_31_0_sva_2 & state_0_2_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_3_sva_1 = plaintext_31_0_sva_3 & state_0_3_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_59_sva_1 = plaintext_63_32_sva_27 & state_0_59_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_4_sva_1 = plaintext_31_0_sva_4 & state_0_4_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_58_sva_1 = plaintext_63_32_sva_26 & state_0_58_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_5_sva_1 = plaintext_31_0_sva_5 & state_0_5_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_57_sva_1 = plaintext_63_32_sva_25 & state_0_57_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_6_sva_1 = plaintext_31_0_sva_6 & state_0_6_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_56_sva_1 = plaintext_63_32_sva_24 & state_0_56_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_7_sva_1 = plaintext_31_0_sva_7 & state_0_7_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_55_sva_1 = plaintext_63_32_sva_23 & state_0_55_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_8_sva_1 = plaintext_31_0_sva_8 & state_0_8_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_54_sva_1 = plaintext_63_32_sva_22 & state_0_54_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_9_sva_1 = plaintext_31_0_sva_9 & state_0_9_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_53_sva_1 = plaintext_63_32_sva_21 & state_0_53_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_52_sva_1 = plaintext_63_32_sva_20 & state_0_52_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_51_sva_1 = plaintext_63_32_sva_19 & state_0_51_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_50_sva_1 = plaintext_63_32_sva_18 & state_0_50_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_49_sva_1 = plaintext_63_32_sva_17 & state_0_49_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_48_sva_1 = plaintext_63_32_sva_16 & state_0_48_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_47_sva_1 = plaintext_63_32_sva_15 & state_0_47_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_46_sva_1 = plaintext_63_32_sva_14 & state_0_46_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_17_sva_1 = plaintext_31_0_sva_17 & state_0_17_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_45_sva_1 = plaintext_63_32_sva_13 & state_0_45_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_44_sva_1 = plaintext_63_32_sva_12 & state_0_44_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_43_sva_1 = plaintext_63_32_sva_11 & state_0_43_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_42_sva_1 = plaintext_63_32_sva_10 & state_0_42_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_41_sva_1 = plaintext_63_32_sva_9 & state_0_41_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_40_sva_1 = plaintext_63_32_sva_8 & state_0_40_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_39_sva_1 = plaintext_63_32_sva_7 & state_0_39_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_38_sva_1 = plaintext_63_32_sva_6 & state_0_38_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_37_sva_1 = plaintext_63_32_sva_5 & state_0_37_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_36_sva_1 = plaintext_63_32_sva_4 & state_0_36_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_35_sva_1 = plaintext_63_32_sva_3 & state_0_35_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_34_sva_1 = plaintext_63_32_sva_2 & state_0_34_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_33_sva_1 = plaintext_63_32_sva_1 & state_0_33_lpi_6;
  assign Encrypt_Top_sbox_and_2_cse_32_sva_1 = plaintext_63_32_sva_0 & state_0_32_lpi_6;
  assign INIT_P12_INIT_P12_xor_8_psp_sva_1 = state_2_0_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0]);
  assign INIT_P12_INIT_P12_xor_7_psp_sva_1 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1]);
  assign INIT_P12_INIT_P12_xor_6_psp_sva_1 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2]);
  assign INIT_P12_INIT_P12_xor_5_psp_sva_1 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3]);
  assign INIT_P12_INIT_P12_xor_4_psp_sva_1 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4]);
  assign INIT_P12_INIT_P12_xor_3_psp_sva_1 = state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5]);
  assign INIT_P12_INIT_P12_xor_2_psp_sva_1 = state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6]);
  assign INIT_P12_INIT_P12_xor_1_psp_sva_1 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7]);
  assign Encrypt_Top_sbox_and_1_cse_63_sva_1 = state_2_63_1_lpi_4 & plaintext_63_32_sva_31;
  assign Encrypt_Top_sbox_and_1_cse_0_sva_1 = INIT_P12_INIT_P12_xor_8_psp_sva_1 &
      plaintext_31_0_sva_0;
  assign Encrypt_Top_sbox_and_1_cse_62_sva_1 = state_2_62_1_lpi_4 & plaintext_63_32_sva_30;
  assign Encrypt_Top_sbox_and_1_cse_1_sva_1 = INIT_P12_INIT_P12_xor_7_psp_sva_1 &
      plaintext_31_0_sva_1;
  assign Encrypt_Top_sbox_and_1_cse_61_sva_1 = state_2_61_1_lpi_4 & plaintext_63_32_sva_29;
  assign Encrypt_Top_sbox_and_1_cse_2_sva_1 = INIT_P12_INIT_P12_xor_6_psp_sva_1 &
      plaintext_31_0_sva_2;
  assign Encrypt_Top_sbox_and_1_cse_60_sva_1 = state_2_60_1_lpi_4 & plaintext_63_32_sva_28;
  assign Encrypt_Top_sbox_and_1_cse_3_sva_1 = INIT_P12_INIT_P12_xor_5_psp_sva_1 &
      plaintext_31_0_sva_3;
  assign Encrypt_Top_sbox_and_1_cse_59_sva_1 = state_2_59_1_lpi_4 & plaintext_63_32_sva_27;
  assign Encrypt_Top_sbox_and_1_cse_4_sva_1 = INIT_P12_INIT_P12_xor_4_psp_sva_1 &
      plaintext_31_0_sva_4;
  assign Encrypt_Top_sbox_and_1_cse_58_sva_1 = state_2_58_1_lpi_4 & plaintext_63_32_sva_26;
  assign Encrypt_Top_sbox_and_1_cse_5_sva_1 = INIT_P12_INIT_P12_xor_3_psp_sva_1 &
      plaintext_31_0_sva_5;
  assign Encrypt_Top_sbox_and_1_cse_57_sva_1 = state_2_57_1_lpi_4 & plaintext_63_32_sva_25;
  assign Encrypt_Top_sbox_and_1_cse_6_sva_1 = INIT_P12_INIT_P12_xor_2_psp_sva_1 &
      plaintext_31_0_sva_6;
  assign Encrypt_Top_sbox_and_1_cse_56_sva_1 = state_2_56_1_lpi_4 & plaintext_63_32_sva_24;
  assign Encrypt_Top_sbox_and_1_cse_7_sva_1 = INIT_P12_INIT_P12_xor_1_psp_sva_1 &
      plaintext_31_0_sva_7;
  assign Encrypt_Top_sbox_and_1_cse_55_sva_1 = state_2_55_1_lpi_4 & plaintext_63_32_sva_23;
  assign Encrypt_Top_sbox_and_1_cse_8_sva_1 = state_2_8_1_lpi_4 & plaintext_31_0_sva_8;
  assign Encrypt_Top_sbox_and_1_cse_54_sva_1 = state_2_54_1_lpi_4 & plaintext_63_32_sva_22;
  assign Encrypt_Top_sbox_and_1_cse_9_sva_1 = state_2_9_1_lpi_4 & plaintext_31_0_sva_9;
  assign Encrypt_Top_sbox_and_1_cse_53_sva_1 = state_2_53_1_lpi_4 & plaintext_63_32_sva_21;
  assign Encrypt_Top_sbox_and_1_cse_10_sva_1 = state_2_10_1_lpi_4 & plaintext_31_0_sva_10;
  assign Encrypt_Top_sbox_and_1_cse_52_sva_1 = state_2_52_1_lpi_4 & plaintext_63_32_sva_20;
  assign Encrypt_Top_sbox_and_1_cse_11_sva_1 = state_2_11_1_lpi_4 & plaintext_31_0_sva_11;
  assign Encrypt_Top_sbox_and_1_cse_51_sva_1 = state_2_51_1_lpi_4 & plaintext_63_32_sva_19;
  assign Encrypt_Top_sbox_and_1_cse_12_sva_1 = state_2_12_1_lpi_4 & plaintext_31_0_sva_12;
  assign Encrypt_Top_sbox_and_1_cse_50_sva_1 = state_2_50_1_lpi_4 & plaintext_63_32_sva_18;
  assign Encrypt_Top_sbox_and_1_cse_13_sva_1 = state_2_13_1_lpi_4 & plaintext_31_0_sva_13;
  assign Encrypt_Top_sbox_and_1_cse_49_sva_1 = state_2_49_1_lpi_4 & plaintext_63_32_sva_17;
  assign Encrypt_Top_sbox_and_1_cse_14_sva_1 = state_2_14_1_lpi_4 & plaintext_31_0_sva_14;
  assign Encrypt_Top_sbox_and_1_cse_48_sva_1 = state_2_48_1_lpi_4 & plaintext_63_32_sva_16;
  assign Encrypt_Top_sbox_and_1_cse_15_sva_1 = state_2_15_1_lpi_4 & plaintext_31_0_sva_15;
  assign Encrypt_Top_sbox_and_1_cse_47_sva_1 = state_2_47_1_lpi_4 & plaintext_63_32_sva_15;
  assign Encrypt_Top_sbox_and_1_cse_16_sva_1 = state_2_16_1_lpi_4 & plaintext_31_0_sva_16;
  assign Encrypt_Top_sbox_and_1_cse_46_sva_1 = state_2_46_1_lpi_4 & plaintext_63_32_sva_14;
  assign Encrypt_Top_sbox_and_1_cse_17_sva_1 = state_2_17_1_lpi_4 & plaintext_31_0_sva_17;
  assign Encrypt_Top_sbox_and_1_cse_45_sva_1 = state_2_45_1_lpi_4 & plaintext_63_32_sva_13;
  assign Encrypt_Top_sbox_and_1_cse_18_sva_1 = state_2_18_1_lpi_4 & plaintext_31_0_sva_18;
  assign Encrypt_Top_sbox_and_1_cse_44_sva_1 = state_2_44_1_lpi_4 & plaintext_63_32_sva_12;
  assign Encrypt_Top_sbox_and_1_cse_19_sva_1 = state_2_19_1_lpi_4 & plaintext_31_0_sva_19;
  assign Encrypt_Top_sbox_and_1_cse_43_sva_1 = state_2_43_1_lpi_4 & plaintext_63_32_sva_11;
  assign Encrypt_Top_sbox_and_1_cse_20_sva_1 = state_2_20_1_lpi_4 & plaintext_31_0_sva_20;
  assign Encrypt_Top_sbox_and_1_cse_42_sva_1 = state_2_42_1_lpi_4 & plaintext_63_32_sva_10;
  assign Encrypt_Top_sbox_and_1_cse_21_sva_1 = state_2_21_1_lpi_4 & plaintext_31_0_sva_21;
  assign Encrypt_Top_sbox_and_1_cse_41_sva_1 = state_2_41_1_lpi_4 & plaintext_63_32_sva_9;
  assign Encrypt_Top_sbox_and_1_cse_22_sva_1 = state_2_22_1_lpi_4 & plaintext_31_0_sva_22;
  assign Encrypt_Top_sbox_and_1_cse_40_sva_1 = state_2_40_1_lpi_4 & plaintext_63_32_sva_8;
  assign Encrypt_Top_sbox_and_1_cse_23_sva_1 = state_2_23_1_lpi_4 & plaintext_31_0_sva_23;
  assign Encrypt_Top_sbox_and_1_cse_39_sva_1 = state_2_39_1_lpi_4 & plaintext_63_32_sva_7;
  assign Encrypt_Top_sbox_and_1_cse_24_sva_1 = state_2_24_1_lpi_4 & plaintext_31_0_sva_24;
  assign Encrypt_Top_sbox_and_1_cse_38_sva_1 = state_2_38_1_lpi_4 & plaintext_63_32_sva_6;
  assign Encrypt_Top_sbox_and_1_cse_25_sva_1 = state_2_25_1_lpi_4 & plaintext_31_0_sva_25;
  assign Encrypt_Top_sbox_and_1_cse_37_sva_1 = state_2_37_1_lpi_4 & plaintext_63_32_sva_5;
  assign Encrypt_Top_sbox_and_1_cse_26_sva_1 = state_2_26_1_lpi_4 & plaintext_31_0_sva_26;
  assign Encrypt_Top_sbox_and_1_cse_36_sva_1 = state_2_36_1_lpi_4 & plaintext_63_32_sva_4;
  assign Encrypt_Top_sbox_and_1_cse_27_sva_1 = state_2_27_1_lpi_4 & plaintext_31_0_sva_27;
  assign Encrypt_Top_sbox_and_1_cse_35_sva_1 = state_2_35_1_lpi_4 & plaintext_63_32_sva_3;
  assign Encrypt_Top_sbox_and_1_cse_28_sva_1 = state_2_28_1_lpi_4 & plaintext_31_0_sva_28;
  assign Encrypt_Top_sbox_and_1_cse_34_sva_1 = state_2_34_1_lpi_4 & plaintext_63_32_sva_2;
  assign Encrypt_Top_sbox_and_1_cse_29_sva_1 = state_2_29_1_lpi_4 & plaintext_31_0_sva_29;
  assign Encrypt_Top_sbox_and_1_cse_33_sva_1 = state_2_33_1_lpi_4 & plaintext_63_32_sva_1;
  assign Encrypt_Top_sbox_and_1_cse_30_sva_1 = state_2_30_1_lpi_4 & plaintext_31_0_sva_30;
  assign Encrypt_Top_sbox_and_1_cse_32_sva_1 = state_2_32_1_lpi_4 & plaintext_63_32_sva_0;
  assign Encrypt_Top_sbox_and_1_cse_31_sva_1 = state_2_31_1_lpi_4 & plaintext_31_0_sva_31;
  assign nl_AD_P6_j_2_0_sva_2 = AD_P6_j_2_0_sva + 3'b001;
  assign AD_P6_j_2_0_sva_2 = nl_AD_P6_j_2_0_sva_2[2:0];
  assign Encrypt_Top_sbox_1_and_cse_62_sva_1 = state_4_4_62_lpi_3 & state_1_1_63_32_lpi_4_30;
  assign Encrypt_Top_sbox_2_and_2_cse_62_sva_1 = state_1_1_63_32_lpi_4_30 & state_0_62_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_61_sva_1 = state_4_4_61_lpi_3 & state_1_1_63_32_lpi_4_29;
  assign Encrypt_Top_sbox_2_and_2_cse_61_sva_1 = state_1_1_63_32_lpi_4_29 & state_0_61_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_60_sva_1 = state_4_4_60_lpi_3 & state_1_1_63_32_lpi_4_28;
  assign Encrypt_Top_sbox_2_and_2_cse_60_sva_1 = state_1_1_63_32_lpi_4_28 & state_0_60_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_59_sva_1 = state_4_4_59_lpi_3 & state_1_1_63_32_lpi_4_27;
  assign Encrypt_Top_sbox_2_and_2_cse_59_sva_1 = state_1_1_63_32_lpi_4_27 & state_0_59_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_10_sva_1 = state_4_4_10_lpi_3 & state_1_1_31_0_lpi_4_10;
  assign Encrypt_Top_sbox_2_and_2_cse_10_sva_1 = state_1_1_31_0_lpi_4_10 & state_0_10_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_11_sva_1 = state_4_4_11_lpi_3 & state_1_1_31_0_lpi_4_11;
  assign Encrypt_Top_sbox_2_and_2_cse_11_sva_1 = state_1_1_31_0_lpi_4_11 & state_0_11_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_12_sva_1 = state_4_4_12_lpi_3 & state_1_1_31_0_lpi_4_12;
  assign Encrypt_Top_sbox_2_and_2_cse_12_sva_1 = state_1_1_31_0_lpi_4_12 & state_0_12_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_13_sva_1 = state_4_4_13_lpi_3 & state_1_1_31_0_lpi_4_13;
  assign Encrypt_Top_sbox_2_and_2_cse_13_sva_1 = state_1_1_31_0_lpi_4_13 & state_0_13_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_14_sva_1 = state_4_4_14_lpi_3 & state_1_1_31_0_lpi_4_14;
  assign Encrypt_Top_sbox_2_and_2_cse_14_sva_1 = state_1_1_31_0_lpi_4_14 & state_0_14_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_15_sva_1 = state_4_4_15_lpi_3 & state_1_1_31_0_lpi_4_15;
  assign Encrypt_Top_sbox_2_and_2_cse_15_sva_1 = state_1_1_31_0_lpi_4_15 & state_0_15_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_16_sva_1 = state_4_4_16_lpi_3 & state_1_1_31_0_lpi_4_16;
  assign Encrypt_Top_sbox_2_and_2_cse_16_sva_1 = state_1_1_31_0_lpi_4_16 & state_0_16_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_17_sva_1 = state_4_4_17_lpi_3 & state_1_1_31_0_lpi_4_17;
  assign Encrypt_Top_sbox_2_and_2_cse_17_sva_1 = state_1_1_31_0_lpi_4_17 & state_0_17_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_18_sva_1 = state_4_4_18_lpi_3 & state_1_1_31_0_lpi_4_18;
  assign Encrypt_Top_sbox_2_and_2_cse_18_sva_1 = state_1_1_31_0_lpi_4_18 & state_0_18_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_44_sva_1 = state_4_4_44_lpi_3 & state_1_1_63_32_lpi_4_12;
  assign Encrypt_Top_sbox_2_and_2_cse_44_sva_1 = state_1_1_63_32_lpi_4_12 & state_0_44_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_19_sva_1 = state_4_4_19_lpi_3 & state_1_1_31_0_lpi_4_19;
  assign Encrypt_Top_sbox_2_and_2_cse_19_sva_1 = state_1_1_31_0_lpi_4_19 & state_0_19_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_20_sva_1 = state_4_4_20_lpi_3 & state_1_1_31_0_lpi_4_20;
  assign Encrypt_Top_sbox_2_and_2_cse_20_sva_1 = state_1_1_31_0_lpi_4_20 & state_0_20_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_42_sva_1 = state_4_4_42_lpi_3 & state_1_1_63_32_lpi_4_10;
  assign Encrypt_Top_sbox_2_and_2_cse_42_sva_1 = state_1_1_63_32_lpi_4_10 & state_0_42_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_21_sva_1 = state_4_4_21_lpi_3 & state_1_1_31_0_lpi_4_21;
  assign Encrypt_Top_sbox_2_and_2_cse_21_sva_1 = state_1_1_31_0_lpi_4_21 & state_0_21_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_41_sva_1 = state_4_4_41_lpi_3 & state_1_1_63_32_lpi_4_9;
  assign Encrypt_Top_sbox_2_and_2_cse_41_sva_1 = state_1_1_63_32_lpi_4_9 & state_0_41_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_22_sva_1 = state_4_4_22_lpi_3 & state_1_1_31_0_lpi_4_22;
  assign Encrypt_Top_sbox_2_and_2_cse_22_sva_1 = state_1_1_31_0_lpi_4_22 & state_0_22_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_23_sva_1 = state_4_4_23_lpi_3 & state_1_1_31_0_lpi_4_23;
  assign Encrypt_Top_sbox_2_and_2_cse_23_sva_1 = state_1_1_31_0_lpi_4_23 & state_0_23_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_24_sva_1 = state_4_4_24_lpi_3 & state_1_1_31_0_lpi_4_24;
  assign Encrypt_Top_sbox_2_and_2_cse_24_sva_1 = state_1_1_31_0_lpi_4_24 & state_0_24_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_25_sva_1 = state_4_4_25_lpi_3 & state_1_1_31_0_lpi_4_25;
  assign Encrypt_Top_sbox_2_and_2_cse_25_sva_1 = state_1_1_31_0_lpi_4_25 & state_0_25_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_26_sva_1 = state_4_4_26_lpi_3 & state_1_1_31_0_lpi_4_26;
  assign Encrypt_Top_sbox_2_and_2_cse_26_sva_1 = state_1_1_31_0_lpi_4_26 & state_0_26_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_27_sva_1 = state_4_4_27_lpi_3 & state_1_1_31_0_lpi_4_27;
  assign Encrypt_Top_sbox_2_and_2_cse_27_sva_1 = state_1_1_31_0_lpi_4_27 & state_0_27_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_28_sva_1 = state_4_4_28_lpi_3 & state_1_1_31_0_lpi_4_28;
  assign Encrypt_Top_sbox_2_and_2_cse_28_sva_1 = state_1_1_31_0_lpi_4_28 & state_0_28_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_29_sva_1 = state_4_4_29_lpi_3 & state_1_1_31_0_lpi_4_29;
  assign Encrypt_Top_sbox_2_and_2_cse_29_sva_1 = state_1_1_31_0_lpi_4_29 & state_0_29_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_30_sva_1 = state_4_4_30_lpi_3 & state_1_1_31_0_lpi_4_30;
  assign Encrypt_Top_sbox_2_and_2_cse_30_sva_1 = state_1_1_31_0_lpi_4_30 & state_0_30_lpi_6;
  assign Encrypt_Top_sbox_1_and_cse_31_sva_1 = state_4_4_31_lpi_3 & state_1_1_31_0_lpi_4_31;
  assign Encrypt_Top_sbox_2_and_2_cse_31_sva_1 = state_1_1_31_0_lpi_4_31 & state_0_31_lpi_6;
  assign AD_P6_AD_P6_xor_8_psp_sva_1 = state_2_0_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]);
  assign AD_P6_AD_P6_xor_7_psp_sva_1 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]);
  assign AD_P6_AD_P6_xor_6_psp_sva_1 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]);
  assign AD_P6_AD_P6_xor_5_psp_sva_1 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]);
  assign AD_P6_AD_P6_xor_4_psp_sva_1 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign AD_P6_AD_P6_xor_3_psp_sva_1 = state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]);
  assign AD_P6_AD_P6_xor_2_psp_sva_1 = state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]);
  assign AD_P6_AD_P6_xor_1_psp_sva_1 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]);
  assign Encrypt_Top_sbox_1_and_1_cse_63_sva_1 = state_2_63_1_lpi_4 & state_1_1_63_32_lpi_4_31;
  assign Encrypt_Top_sbox_1_and_1_cse_0_sva_1 = AD_P6_AD_P6_xor_8_psp_sva_1 & state_1_1_31_0_lpi_4_0;
  assign Encrypt_Top_sbox_1_and_1_cse_62_sva_1 = state_2_62_1_lpi_4 & state_1_1_63_32_lpi_4_30;
  assign Encrypt_Top_sbox_1_and_1_cse_1_sva_1 = AD_P6_AD_P6_xor_7_psp_sva_1 & state_1_1_31_0_lpi_4_1;
  assign Encrypt_Top_sbox_1_and_1_cse_61_sva_1 = state_2_61_1_lpi_4 & state_1_1_63_32_lpi_4_29;
  assign Encrypt_Top_sbox_1_and_1_cse_2_sva_1 = AD_P6_AD_P6_xor_6_psp_sva_1 & state_1_1_31_0_lpi_4_2;
  assign Encrypt_Top_sbox_1_and_1_cse_60_sva_1 = state_2_60_1_lpi_4 & state_1_1_63_32_lpi_4_28;
  assign Encrypt_Top_sbox_1_and_1_cse_3_sva_1 = AD_P6_AD_P6_xor_5_psp_sva_1 & state_1_1_31_0_lpi_4_3;
  assign Encrypt_Top_sbox_1_and_1_cse_59_sva_1 = state_2_59_1_lpi_4 & state_1_1_63_32_lpi_4_27;
  assign Encrypt_Top_sbox_1_and_1_cse_4_sva_1 = AD_P6_AD_P6_xor_4_psp_sva_1 & state_1_1_31_0_lpi_4_4;
  assign Encrypt_Top_sbox_1_and_1_cse_58_sva_1 = state_2_58_1_lpi_4 & state_1_1_63_32_lpi_4_26;
  assign Encrypt_Top_sbox_1_and_1_cse_5_sva_1 = AD_P6_AD_P6_xor_3_psp_sva_1 & state_1_1_31_0_lpi_4_5;
  assign Encrypt_Top_sbox_1_and_1_cse_57_sva_1 = state_2_57_1_lpi_4 & state_1_1_63_32_lpi_4_25;
  assign Encrypt_Top_sbox_1_and_1_cse_6_sva_1 = AD_P6_AD_P6_xor_2_psp_sva_1 & state_1_1_31_0_lpi_4_6;
  assign Encrypt_Top_sbox_1_and_1_cse_56_sva_1 = state_2_56_1_lpi_4 & state_1_1_63_32_lpi_4_24;
  assign Encrypt_Top_sbox_1_and_1_cse_7_sva_1 = AD_P6_AD_P6_xor_1_psp_sva_1 & state_1_1_31_0_lpi_4_7;
  assign Encrypt_Top_sbox_1_and_1_cse_55_sva_1 = state_2_55_1_lpi_4 & state_1_1_63_32_lpi_4_23;
  assign Encrypt_Top_sbox_1_and_1_cse_8_sva_1 = state_2_8_1_lpi_4 & state_1_1_31_0_lpi_4_8;
  assign Encrypt_Top_sbox_1_and_1_cse_54_sva_1 = state_2_54_1_lpi_4 & state_1_1_63_32_lpi_4_22;
  assign Encrypt_Top_sbox_1_and_1_cse_9_sva_1 = state_2_9_1_lpi_4 & state_1_1_31_0_lpi_4_9;
  assign Encrypt_Top_sbox_1_and_1_cse_53_sva_1 = state_2_53_1_lpi_4 & state_1_1_63_32_lpi_4_21;
  assign Encrypt_Top_sbox_1_and_1_cse_10_sva_1 = state_2_10_1_lpi_4 & state_1_1_31_0_lpi_4_10;
  assign Encrypt_Top_sbox_1_and_1_cse_52_sva_1 = state_2_52_1_lpi_4 & state_1_1_63_32_lpi_4_20;
  assign Encrypt_Top_sbox_1_and_1_cse_11_sva_1 = state_2_11_1_lpi_4 & state_1_1_31_0_lpi_4_11;
  assign Encrypt_Top_sbox_1_and_1_cse_51_sva_1 = state_2_51_1_lpi_4 & state_1_1_63_32_lpi_4_19;
  assign Encrypt_Top_sbox_1_and_1_cse_12_sva_1 = state_2_12_1_lpi_4 & state_1_1_31_0_lpi_4_12;
  assign Encrypt_Top_sbox_1_and_1_cse_50_sva_1 = state_2_50_1_lpi_4 & state_1_1_63_32_lpi_4_18;
  assign Encrypt_Top_sbox_1_and_1_cse_13_sva_1 = state_2_13_1_lpi_4 & state_1_1_31_0_lpi_4_13;
  assign Encrypt_Top_sbox_1_and_1_cse_49_sva_1 = state_2_49_1_lpi_4 & state_1_1_63_32_lpi_4_17;
  assign Encrypt_Top_sbox_1_and_1_cse_14_sva_1 = state_2_14_1_lpi_4 & state_1_1_31_0_lpi_4_14;
  assign Encrypt_Top_sbox_1_and_1_cse_48_sva_1 = state_2_48_1_lpi_4 & state_1_1_63_32_lpi_4_16;
  assign Encrypt_Top_sbox_1_and_1_cse_15_sva_1 = state_2_15_1_lpi_4 & state_1_1_31_0_lpi_4_15;
  assign Encrypt_Top_sbox_1_and_1_cse_47_sva_1 = state_2_47_1_lpi_4 & state_1_1_63_32_lpi_4_15;
  assign Encrypt_Top_sbox_1_and_1_cse_16_sva_1 = state_2_16_1_lpi_4 & state_1_1_31_0_lpi_4_16;
  assign Encrypt_Top_sbox_1_and_1_cse_46_sva_1 = state_2_46_1_lpi_4 & state_1_1_63_32_lpi_4_14;
  assign Encrypt_Top_sbox_1_and_1_cse_17_sva_1 = state_2_17_1_lpi_4 & state_1_1_31_0_lpi_4_17;
  assign Encrypt_Top_sbox_1_and_1_cse_45_sva_1 = state_2_45_1_lpi_4 & state_1_1_63_32_lpi_4_13;
  assign Encrypt_Top_sbox_1_and_1_cse_18_sva_1 = state_2_18_1_lpi_4 & state_1_1_31_0_lpi_4_18;
  assign Encrypt_Top_sbox_1_and_1_cse_44_sva_1 = state_2_44_1_lpi_4 & state_1_1_63_32_lpi_4_12;
  assign Encrypt_Top_sbox_1_and_1_cse_19_sva_1 = state_2_19_1_lpi_4 & state_1_1_31_0_lpi_4_19;
  assign Encrypt_Top_sbox_1_and_1_cse_43_sva_1 = state_2_43_1_lpi_4 & state_1_1_63_32_lpi_4_11;
  assign Encrypt_Top_sbox_1_and_1_cse_20_sva_1 = state_2_20_1_lpi_4 & state_1_1_31_0_lpi_4_20;
  assign Encrypt_Top_sbox_1_and_1_cse_42_sva_1 = state_2_42_1_lpi_4 & state_1_1_63_32_lpi_4_10;
  assign Encrypt_Top_sbox_1_and_1_cse_21_sva_1 = state_2_21_1_lpi_4 & state_1_1_31_0_lpi_4_21;
  assign Encrypt_Top_sbox_1_and_1_cse_41_sva_1 = state_2_41_1_lpi_4 & state_1_1_63_32_lpi_4_9;
  assign Encrypt_Top_sbox_1_and_1_cse_22_sva_1 = state_2_22_1_lpi_4 & state_1_1_31_0_lpi_4_22;
  assign Encrypt_Top_sbox_1_and_1_cse_40_sva_1 = state_2_40_1_lpi_4 & state_1_1_63_32_lpi_4_8;
  assign Encrypt_Top_sbox_1_and_1_cse_23_sva_1 = state_2_23_1_lpi_4 & state_1_1_31_0_lpi_4_23;
  assign Encrypt_Top_sbox_1_and_1_cse_39_sva_1 = state_2_39_1_lpi_4 & state_1_1_63_32_lpi_4_7;
  assign Encrypt_Top_sbox_1_and_1_cse_24_sva_1 = state_2_24_1_lpi_4 & state_1_1_31_0_lpi_4_24;
  assign Encrypt_Top_sbox_1_and_1_cse_38_sva_1 = state_2_38_1_lpi_4 & state_1_1_63_32_lpi_4_6;
  assign Encrypt_Top_sbox_1_and_1_cse_25_sva_1 = state_2_25_1_lpi_4 & state_1_1_31_0_lpi_4_25;
  assign Encrypt_Top_sbox_1_and_1_cse_37_sva_1 = state_2_37_1_lpi_4 & state_1_1_63_32_lpi_4_5;
  assign Encrypt_Top_sbox_1_and_1_cse_26_sva_1 = state_2_26_1_lpi_4 & state_1_1_31_0_lpi_4_26;
  assign Encrypt_Top_sbox_1_and_1_cse_36_sva_1 = state_2_36_1_lpi_4 & state_1_1_63_32_lpi_4_4;
  assign Encrypt_Top_sbox_1_and_1_cse_27_sva_1 = state_2_27_1_lpi_4 & state_1_1_31_0_lpi_4_27;
  assign Encrypt_Top_sbox_1_and_1_cse_35_sva_1 = state_2_35_1_lpi_4 & state_1_1_63_32_lpi_4_3;
  assign Encrypt_Top_sbox_1_and_1_cse_28_sva_1 = state_2_28_1_lpi_4 & state_1_1_31_0_lpi_4_28;
  assign Encrypt_Top_sbox_1_and_1_cse_34_sva_1 = state_2_34_1_lpi_4 & state_1_1_63_32_lpi_4_2;
  assign Encrypt_Top_sbox_1_and_1_cse_29_sva_1 = state_2_29_1_lpi_4 & state_1_1_31_0_lpi_4_29;
  assign Encrypt_Top_sbox_1_and_1_cse_33_sva_1 = state_2_33_1_lpi_4 & state_1_1_63_32_lpi_4_1;
  assign Encrypt_Top_sbox_1_and_1_cse_30_sva_1 = state_2_30_1_lpi_4 & state_1_1_31_0_lpi_4_30;
  assign Encrypt_Top_sbox_1_and_1_cse_32_sva_1 = state_2_32_1_lpi_4 & state_1_1_63_32_lpi_4_0;
  assign Encrypt_Top_sbox_1_and_1_cse_31_sva_1 = state_2_31_1_lpi_4 & state_1_1_31_0_lpi_4_31;
  assign ENC_P6_ENC_P6_xor_8_psp_sva_1 = state_2_0_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]);
  assign ENC_P6_ENC_P6_xor_7_psp_sva_1 = state_2_1_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]);
  assign ENC_P6_ENC_P6_xor_6_psp_sva_1 = state_2_2_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]);
  assign ENC_P6_ENC_P6_xor_5_psp_sva_1 = state_2_3_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]);
  assign ENC_P6_ENC_P6_xor_4_psp_sva_1 = state_2_4_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign ENC_P6_ENC_P6_xor_3_psp_sva_1 = state_2_5_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]);
  assign ENC_P6_ENC_P6_xor_2_psp_sva_1 = state_2_6_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]);
  assign ENC_P6_ENC_P6_xor_1_psp_sva_1 = state_2_7_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]);
  assign Encrypt_Top_sbox_2_and_1_cse_0_sva_1 = ENC_P6_ENC_P6_xor_8_psp_sva_1 & state_1_1_31_0_lpi_4_0;
  assign Encrypt_Top_sbox_2_and_1_cse_1_sva_1 = ENC_P6_ENC_P6_xor_7_psp_sva_1 & state_1_1_31_0_lpi_4_1;
  assign Encrypt_Top_sbox_2_and_1_cse_2_sva_1 = ENC_P6_ENC_P6_xor_6_psp_sva_1 & state_1_1_31_0_lpi_4_2;
  assign Encrypt_Top_sbox_2_and_1_cse_3_sva_1 = ENC_P6_ENC_P6_xor_5_psp_sva_1 & state_1_1_31_0_lpi_4_3;
  assign Encrypt_Top_sbox_2_and_1_cse_4_sva_1 = ENC_P6_ENC_P6_xor_4_psp_sva_1 & state_1_1_31_0_lpi_4_4;
  assign Encrypt_Top_sbox_2_and_1_cse_5_sva_1 = ENC_P6_ENC_P6_xor_3_psp_sva_1 & state_1_1_31_0_lpi_4_5;
  assign Encrypt_Top_sbox_2_and_1_cse_6_sva_1 = ENC_P6_ENC_P6_xor_2_psp_sva_1 & state_1_1_31_0_lpi_4_6;
  assign Encrypt_Top_sbox_2_and_1_cse_7_sva_1 = ENC_P6_ENC_P6_xor_1_psp_sva_1 & state_1_1_31_0_lpi_4_7;
  assign Encrypt_Top_sbox_3_and_cse_50_sva_1 = state_4_4_50_lpi_3 & state_1_1_63_32_lpi_4_23;
  assign Encrypt_Top_sbox_3_and_2_cse_50_sva_1 = state_1_1_63_32_lpi_4_23 & state_0_50_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_48_sva_1 = state_4_4_48_lpi_3 & state_1_1_63_32_lpi_4_21;
  assign Encrypt_Top_sbox_3_and_2_cse_48_sva_1 = state_1_1_63_32_lpi_4_21 & state_0_48_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_47_sva_1 = state_4_4_47_lpi_3 & state_1_1_63_32_lpi_4_20;
  assign Encrypt_Top_sbox_3_and_2_cse_47_sva_1 = state_1_1_63_32_lpi_4_20 & state_0_47_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_45_sva_1 = state_4_4_45_lpi_3 & state_1_1_63_32_lpi_4_19;
  assign Encrypt_Top_sbox_3_and_2_cse_45_sva_1 = state_1_1_63_32_lpi_4_19 & state_0_45_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_43_sva_1 = state_4_4_43_lpi_3 & state_1_1_63_32_lpi_4_17;
  assign Encrypt_Top_sbox_3_and_2_cse_43_sva_1 = state_1_1_63_32_lpi_4_17 & state_0_43_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_41_sva_1 = state_4_4_41_lpi_3 & state_1_1_63_32_lpi_4_15;
  assign Encrypt_Top_sbox_3_and_2_cse_41_sva_1 = state_1_1_63_32_lpi_4_15 & state_0_41_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_39_sva_1 = state_4_4_39_lpi_3 & state_1_1_63_32_lpi_4_13;
  assign Encrypt_Top_sbox_3_and_2_cse_39_sva_1 = state_1_1_63_32_lpi_4_13 & state_0_39_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_37_sva_1 = state_4_4_37_lpi_3 & state_1_1_63_32_lpi_4_11;
  assign Encrypt_Top_sbox_3_and_2_cse_37_sva_1 = state_1_1_63_32_lpi_4_11 & state_0_37_lpi_6;
  assign Encrypt_Top_sbox_3_and_cse_36_sva_1 = state_4_4_36_lpi_3 & state_1_1_63_32_lpi_4_10;
  assign Encrypt_Top_sbox_3_and_2_cse_36_sva_1 = state_1_1_63_32_lpi_4_10 & state_0_36_lpi_6;
  assign Encrypt_Top_sbox_3_and_1_cse_32_sva_1 = state_2_32_1_lpi_4 & state_1_1_31_0_lpi_4_8;
  assign Encrypt_Top_sbox_3_and_1_cse_33_sva_1 = state_2_33_1_lpi_4 & state_1_1_31_0_lpi_4_9;
  assign Encrypt_Top_sbox_3_and_1_cse_34_sva_1 = state_2_34_1_lpi_4 & state_1_1_63_32_lpi_4_0;
  assign Encrypt_Top_sbox_3_and_1_cse_35_sva_1 = state_2_35_1_lpi_4 & state_1_1_63_32_lpi_4_1;
  assign Encrypt_Top_sbox_3_and_1_cse_36_sva_1 = state_2_36_1_lpi_4 & state_1_1_63_32_lpi_4_10;
  assign Encrypt_Top_sbox_3_and_1_cse_37_sva_1 = state_2_37_1_lpi_4 & state_1_1_63_32_lpi_4_11;
  assign Encrypt_Top_sbox_3_and_1_cse_38_sva_1 = state_2_38_1_lpi_4 & state_1_1_63_32_lpi_4_12;
  assign Encrypt_Top_sbox_3_and_1_cse_39_sva_1 = state_2_39_1_lpi_4 & state_1_1_63_32_lpi_4_13;
  assign Encrypt_Top_sbox_3_and_1_cse_40_sva_1 = state_2_40_1_lpi_4 & state_1_1_63_32_lpi_4_14;
  assign Encrypt_Top_sbox_3_and_1_cse_41_sva_1 = state_2_41_1_lpi_4 & state_1_1_63_32_lpi_4_15;
  assign Encrypt_Top_sbox_3_and_1_cse_42_sva_1 = state_2_42_1_lpi_4 & state_1_1_63_32_lpi_4_16;
  assign Encrypt_Top_sbox_3_and_1_cse_43_sva_1 = state_2_43_1_lpi_4 & state_1_1_63_32_lpi_4_17;
  assign Encrypt_Top_sbox_3_and_1_cse_44_sva_1 = state_2_44_1_lpi_4 & state_1_1_63_32_lpi_4_18;
  assign Encrypt_Top_sbox_3_and_1_cse_45_sva_1 = state_2_45_1_lpi_4 & state_1_1_63_32_lpi_4_19;
  assign Encrypt_Top_sbox_3_and_1_cse_46_sva_1 = state_2_46_1_lpi_4 & state_1_1_63_32_lpi_4_2;
  assign Encrypt_Top_sbox_3_and_1_cse_47_sva_1 = state_2_47_1_lpi_4 & state_1_1_63_32_lpi_4_20;
  assign Encrypt_Top_sbox_3_and_1_cse_48_sva_1 = state_2_48_1_lpi_4 & state_1_1_63_32_lpi_4_21;
  assign Encrypt_Top_sbox_3_and_1_cse_49_sva_1 = state_2_49_1_lpi_4 & state_1_1_63_32_lpi_4_22;
  assign Encrypt_Top_sbox_3_and_1_cse_50_sva_1 = state_2_50_1_lpi_4 & state_1_1_63_32_lpi_4_23;
  assign Encrypt_Top_sbox_3_and_1_cse_51_sva_1 = state_2_51_1_lpi_4 & state_1_1_63_32_lpi_4_24;
  assign Encrypt_Top_sbox_3_and_1_cse_52_sva_1 = state_2_52_1_lpi_4 & state_1_1_63_32_lpi_4_25;
  assign Encrypt_Top_sbox_3_and_1_cse_53_sva_1 = state_2_53_1_lpi_4 & state_1_1_63_32_lpi_4_26;
  assign Encrypt_Top_sbox_3_and_1_cse_9_sva_1 = state_2_9_1_lpi_4 & state_1_1_63_32_lpi_4_9;
  assign Encrypt_Top_sbox_3_and_1_cse_54_sva_1 = state_2_54_1_lpi_4 & state_1_1_63_32_lpi_4_27;
  assign Encrypt_Top_sbox_3_and_1_cse_8_sva_1 = state_2_8_1_lpi_4 & state_1_1_63_32_lpi_4_8;
  assign Encrypt_Top_sbox_3_and_1_cse_55_sva_1 = state_2_55_1_lpi_4 & state_1_1_63_32_lpi_4_28;
  assign Encrypt_Top_sbox_3_and_1_cse_7_sva_1 = INIT_P12_INIT_P12_xor_1_psp_sva_1
      & state_1_1_31_0_lpi_4_7;
  assign Encrypt_Top_sbox_3_and_1_cse_56_sva_1 = state_2_56_1_lpi_4 & state_1_1_63_32_lpi_4_29;
  assign Encrypt_Top_sbox_3_and_1_cse_6_sva_1 = INIT_P12_INIT_P12_xor_2_psp_sva_1
      & state_1_1_31_0_lpi_4_6;
  assign Encrypt_Top_sbox_3_and_1_cse_57_sva_1 = state_2_57_1_lpi_4 & state_1_1_63_32_lpi_4_3;
  assign Encrypt_Top_sbox_3_and_1_cse_5_sva_1 = INIT_P12_INIT_P12_xor_3_psp_sva_1
      & state_1_1_31_0_lpi_4_5;
  assign Encrypt_Top_sbox_3_and_1_cse_58_sva_1 = state_2_58_1_lpi_4 & state_1_1_63_32_lpi_4_30;
  assign Encrypt_Top_sbox_3_and_1_cse_4_sva_1 = INIT_P12_INIT_P12_xor_4_psp_sva_1
      & state_1_1_31_0_lpi_4_4;
  assign Encrypt_Top_sbox_3_and_1_cse_59_sva_1 = state_2_59_1_lpi_4 & state_1_1_63_32_lpi_4_31;
  assign Encrypt_Top_sbox_3_and_1_cse_3_sva_1 = INIT_P12_INIT_P12_xor_5_psp_sva_1
      & state_1_1_31_0_lpi_4_3;
  assign Encrypt_Top_sbox_3_and_1_cse_60_sva_1 = state_2_60_1_lpi_4 & state_1_1_63_32_lpi_4_4;
  assign Encrypt_Top_sbox_3_and_1_cse_2_sva_1 = INIT_P12_INIT_P12_xor_6_psp_sva_1
      & state_1_1_31_0_lpi_4_2;
  assign Encrypt_Top_sbox_3_and_1_cse_61_sva_1 = state_2_61_1_lpi_4 & state_1_1_63_32_lpi_4_5;
  assign Encrypt_Top_sbox_3_and_1_cse_1_sva_1 = INIT_P12_INIT_P12_xor_7_psp_sva_1
      & state_1_1_31_0_lpi_4_1;
  assign Encrypt_Top_sbox_3_and_1_cse_62_sva_1 = state_2_62_1_lpi_4 & state_1_1_63_32_lpi_4_6;
  assign Encrypt_Top_sbox_3_and_1_cse_0_sva_1 = INIT_P12_INIT_P12_xor_8_psp_sva_1
      & state_1_1_31_0_lpi_4_0;
  assign Encrypt_Top_sbox_3_and_1_cse_63_sva_1 = state_2_63_1_lpi_4 & state_1_1_63_32_lpi_4_7;
  assign Encrypt_Top_sbox_2_and_516 = state_4_4_63_lpi_3 & state_0_63_lpi_6;
  assign Encrypt_Top_sbox_2_and_518 = state_3_63_lpi_3 & state_0_63_lpi_6;
  assign Encrypt_Top_sbox_1_and_516 = state_2_63_1_lpi_4 & state_3_63_lpi_3;
  assign Encrypt_Top_sbox_2_and_520 = state_4_4_0_lpi_3 & state_0_0_lpi_6;
  assign Encrypt_Top_sbox_2_and_522 = state_3_0_lpi_3 & state_0_0_lpi_6;
  assign Encrypt_Top_sbox_2_and_524 = state_4_4_62_lpi_3 & state_0_62_lpi_6;
  assign Encrypt_Top_sbox_2_and_526 = state_3_62_lpi_3 & state_0_62_lpi_6;
  assign Encrypt_Top_sbox_1_and_518 = state_2_62_1_lpi_4 & state_3_62_lpi_3;
  assign Encrypt_Top_sbox_2_and_528 = state_4_4_1_lpi_3 & state_0_1_lpi_6;
  assign Encrypt_Top_sbox_2_and_530 = state_3_1_lpi_3 & state_0_1_lpi_6;
  assign Encrypt_Top_sbox_2_and_532 = state_4_4_61_lpi_3 & state_0_61_lpi_6;
  assign Encrypt_Top_sbox_2_and_534 = state_3_61_lpi_3 & state_0_61_lpi_6;
  assign Encrypt_Top_sbox_1_and_520 = state_2_61_1_lpi_4 & state_3_61_lpi_3;
  assign Encrypt_Top_sbox_2_and_536 = state_4_4_2_lpi_3 & state_0_2_lpi_6;
  assign Encrypt_Top_sbox_2_and_538 = state_3_2_lpi_3 & state_0_2_lpi_6;
  assign Encrypt_Top_sbox_2_and_540 = state_4_4_60_lpi_3 & state_0_60_lpi_6;
  assign Encrypt_Top_sbox_2_and_542 = state_3_60_lpi_3 & state_0_60_lpi_6;
  assign Encrypt_Top_sbox_1_and_522 = state_2_60_1_lpi_4 & state_3_60_lpi_3;
  assign Encrypt_Top_sbox_2_and_544 = state_4_4_3_lpi_3 & state_0_3_lpi_6;
  assign Encrypt_Top_sbox_2_and_546 = state_3_3_lpi_3 & state_0_3_lpi_6;
  assign Encrypt_Top_sbox_2_and_548 = state_4_4_59_lpi_3 & state_0_59_lpi_6;
  assign Encrypt_Top_sbox_2_and_550 = state_3_59_lpi_3 & state_0_59_lpi_6;
  assign Encrypt_Top_sbox_1_and_524 = state_2_59_1_lpi_4 & state_3_59_lpi_3;
  assign Encrypt_Top_sbox_2_and_552 = state_4_4_4_lpi_3 & state_0_4_lpi_6;
  assign Encrypt_Top_sbox_2_and_554 = state_3_4_lpi_3 & state_0_4_lpi_6;
  assign Encrypt_Top_sbox_2_and_556 = state_4_4_58_lpi_3 & state_0_58_lpi_6;
  assign Encrypt_Top_sbox_2_and_558 = state_3_58_lpi_3 & state_0_58_lpi_6;
  assign Encrypt_Top_sbox_1_and_526 = state_2_58_1_lpi_4 & state_3_58_lpi_3;
  assign Encrypt_Top_sbox_2_and_560 = state_4_4_5_lpi_3 & state_0_5_lpi_6;
  assign Encrypt_Top_sbox_2_and_562 = state_3_5_lpi_3 & state_0_5_lpi_6;
  assign Encrypt_Top_sbox_2_and_564 = state_4_4_57_lpi_3 & state_0_57_lpi_6;
  assign Encrypt_Top_sbox_2_and_566 = state_3_57_lpi_3 & state_0_57_lpi_6;
  assign Encrypt_Top_sbox_1_and_528 = state_2_57_1_lpi_4 & state_3_57_lpi_3;
  assign Encrypt_Top_sbox_2_and_568 = state_4_4_6_lpi_3 & state_0_6_lpi_6;
  assign Encrypt_Top_sbox_2_and_570 = state_3_6_lpi_3 & state_0_6_lpi_6;
  assign Encrypt_Top_sbox_2_and_572 = state_4_4_56_lpi_3 & state_0_56_lpi_6;
  assign Encrypt_Top_sbox_2_and_574 = state_3_56_lpi_3 & state_0_56_lpi_6;
  assign Encrypt_Top_sbox_1_and_530 = state_2_56_1_lpi_4 & state_3_56_lpi_3;
  assign Encrypt_Top_sbox_2_and_576 = state_4_4_7_lpi_3 & state_0_7_lpi_6;
  assign Encrypt_Top_sbox_2_and_578 = state_3_7_lpi_3 & state_0_7_lpi_6;
  assign Encrypt_Top_sbox_2_and_580 = state_4_4_55_lpi_3 & state_0_55_lpi_6;
  assign Encrypt_Top_sbox_2_and_582 = state_3_55_lpi_3 & state_0_55_lpi_6;
  assign Encrypt_Top_sbox_1_and_532 = state_2_55_1_lpi_4 & state_3_55_lpi_3;
  assign Encrypt_Top_sbox_2_and_584 = state_4_4_8_lpi_3 & state_0_8_lpi_6;
  assign Encrypt_Top_sbox_2_and_586 = state_3_8_lpi_3 & state_0_8_lpi_6;
  assign Encrypt_Top_sbox_1_and_534 = state_2_8_1_lpi_4 & state_3_8_lpi_3;
  assign Encrypt_Top_sbox_2_and_588 = state_4_4_54_lpi_3 & state_0_54_lpi_6;
  assign Encrypt_Top_sbox_2_and_590 = state_3_54_lpi_3 & state_0_54_lpi_6;
  assign Encrypt_Top_sbox_1_and_536 = state_2_54_1_lpi_4 & state_3_54_lpi_3;
  assign Encrypt_Top_sbox_2_and_592 = state_4_4_9_lpi_3 & state_0_9_lpi_6;
  assign Encrypt_Top_sbox_2_and_594 = state_3_9_lpi_3 & state_0_9_lpi_6;
  assign Encrypt_Top_sbox_1_and_538 = state_2_9_1_lpi_4 & state_3_9_lpi_3;
  assign Encrypt_Top_sbox_2_and_596 = state_4_4_53_lpi_3 & state_0_53_lpi_6;
  assign Encrypt_Top_sbox_2_and_598 = state_3_53_lpi_3 & state_0_53_lpi_6;
  assign Encrypt_Top_sbox_1_and_540 = state_2_53_1_lpi_4 & state_3_53_lpi_3;
  assign Encrypt_Top_sbox_2_and_600 = state_4_4_10_lpi_3 & state_0_10_lpi_6;
  assign Encrypt_Top_sbox_2_and_602 = state_3_10_lpi_3 & state_0_10_lpi_6;
  assign Encrypt_Top_sbox_2_and_604 = state_4_4_52_lpi_3 & state_0_52_lpi_6;
  assign Encrypt_Top_sbox_2_and_606 = state_3_52_lpi_3 & state_0_52_lpi_6;
  assign Encrypt_Top_sbox_1_and_544 = state_2_52_1_lpi_4 & state_3_52_lpi_3;
  assign Encrypt_Top_sbox_2_and_608 = state_4_4_11_lpi_3 & state_0_11_lpi_6;
  assign Encrypt_Top_sbox_2_and_610 = state_3_11_lpi_3 & state_0_11_lpi_6;
  assign Encrypt_Top_sbox_2_and_612 = state_4_4_51_lpi_3 & state_0_51_lpi_6;
  assign Encrypt_Top_sbox_2_and_614 = state_3_51_lpi_3 & state_0_51_lpi_6;
  assign Encrypt_Top_sbox_1_and_548 = state_2_51_1_lpi_4 & state_3_51_lpi_3;
  assign Encrypt_Top_sbox_2_and_616 = state_4_4_12_lpi_3 & state_0_12_lpi_6;
  assign Encrypt_Top_sbox_2_and_618 = state_3_12_lpi_3 & state_0_12_lpi_6;
  assign Encrypt_Top_sbox_2_and_620 = state_4_4_50_lpi_3 & state_0_50_lpi_6;
  assign Encrypt_Top_sbox_2_and_622 = state_3_50_lpi_3 & state_0_50_lpi_6;
  assign Encrypt_Top_sbox_1_and_552 = state_2_50_1_lpi_4 & state_3_50_lpi_3;
  assign Encrypt_Top_sbox_2_and_624 = state_4_4_13_lpi_3 & state_0_13_lpi_6;
  assign Encrypt_Top_sbox_2_and_626 = state_3_13_lpi_3 & state_0_13_lpi_6;
  assign Encrypt_Top_sbox_2_and_628 = state_4_4_49_lpi_3 & state_0_49_lpi_6;
  assign Encrypt_Top_sbox_2_and_630 = state_3_49_lpi_3 & state_0_49_lpi_6;
  assign Encrypt_Top_sbox_1_and_556 = state_2_49_1_lpi_4 & state_3_49_lpi_3;
  assign Encrypt_Top_sbox_2_and_632 = state_4_4_14_lpi_3 & state_0_14_lpi_6;
  assign Encrypt_Top_sbox_2_and_634 = state_3_14_lpi_3 & state_0_14_lpi_6;
  assign Encrypt_Top_sbox_2_and_636 = state_4_4_48_lpi_3 & state_0_48_lpi_6;
  assign Encrypt_Top_sbox_2_and_638 = state_3_48_lpi_3 & state_0_48_lpi_6;
  assign Encrypt_Top_sbox_1_and_560 = state_2_48_1_lpi_4 & state_3_48_lpi_3;
  assign Encrypt_Top_sbox_2_and_640 = state_4_4_15_lpi_3 & state_0_15_lpi_6;
  assign Encrypt_Top_sbox_2_and_642 = state_3_15_lpi_3 & state_0_15_lpi_6;
  assign Encrypt_Top_sbox_2_and_644 = state_4_4_47_lpi_3 & state_0_47_lpi_6;
  assign Encrypt_Top_sbox_2_and_646 = state_3_47_lpi_3 & state_0_47_lpi_6;
  assign Encrypt_Top_sbox_1_and_564 = state_2_47_1_lpi_4 & state_3_47_lpi_3;
  assign Encrypt_Top_sbox_2_and_648 = state_4_4_16_lpi_3 & state_0_16_lpi_6;
  assign Encrypt_Top_sbox_2_and_650 = state_3_16_lpi_3 & state_0_16_lpi_6;
  assign Encrypt_Top_sbox_2_and_652 = state_4_4_46_lpi_3 & state_0_46_lpi_6;
  assign Encrypt_Top_sbox_2_and_654 = state_3_46_lpi_3 & state_0_46_lpi_6;
  assign Encrypt_Top_sbox_1_and_568 = state_2_46_1_lpi_4 & state_3_46_lpi_3;
  assign Encrypt_Top_sbox_2_and_656 = state_4_4_17_lpi_3 & state_0_17_lpi_6;
  assign Encrypt_Top_sbox_2_and_658 = state_3_17_lpi_3 & state_0_17_lpi_6;
  assign Encrypt_Top_sbox_2_and_660 = state_4_4_45_lpi_3 & state_0_45_lpi_6;
  assign Encrypt_Top_sbox_2_and_662 = state_3_45_lpi_3 & state_0_45_lpi_6;
  assign Encrypt_Top_sbox_1_and_572 = state_2_45_1_lpi_4 & state_3_45_lpi_3;
  assign Encrypt_Top_sbox_2_and_664 = state_4_4_18_lpi_3 & state_0_18_lpi_6;
  assign Encrypt_Top_sbox_2_and_666 = state_3_18_lpi_3 & state_0_18_lpi_6;
  assign Encrypt_Top_sbox_2_and_668 = state_4_4_44_lpi_3 & state_0_44_lpi_6;
  assign Encrypt_Top_sbox_2_and_670 = state_3_44_lpi_3 & state_0_44_lpi_6;
  assign Encrypt_Top_sbox_1_and_576 = state_2_44_1_lpi_4 & state_3_44_lpi_3;
  assign Encrypt_Top_sbox_2_and_672 = state_4_4_19_lpi_3 & state_0_19_lpi_6;
  assign Encrypt_Top_sbox_2_and_674 = state_3_19_lpi_3 & state_0_19_lpi_6;
  assign Encrypt_Top_sbox_2_and_676 = state_4_4_43_lpi_3 & state_0_43_lpi_6;
  assign Encrypt_Top_sbox_2_and_678 = state_3_43_lpi_3 & state_0_43_lpi_6;
  assign Encrypt_Top_sbox_1_and_580 = state_2_43_1_lpi_4 & state_3_43_lpi_3;
  assign Encrypt_Top_sbox_2_and_680 = state_4_4_20_lpi_3 & state_0_20_lpi_6;
  assign Encrypt_Top_sbox_2_and_682 = state_3_20_lpi_3 & state_0_20_lpi_6;
  assign Encrypt_Top_sbox_2_and_684 = state_4_4_42_lpi_3 & state_0_42_lpi_6;
  assign Encrypt_Top_sbox_2_and_686 = state_3_42_lpi_3 & state_0_42_lpi_6;
  assign Encrypt_Top_sbox_1_and_584 = state_2_42_1_lpi_4 & state_3_42_lpi_3;
  assign Encrypt_Top_sbox_2_and_688 = state_4_4_21_lpi_3 & state_0_21_lpi_6;
  assign Encrypt_Top_sbox_2_and_690 = state_3_21_lpi_3 & state_0_21_lpi_6;
  assign Encrypt_Top_sbox_2_and_692 = state_4_4_41_lpi_3 & state_0_41_lpi_6;
  assign Encrypt_Top_sbox_2_and_694 = state_3_41_lpi_3 & state_0_41_lpi_6;
  assign Encrypt_Top_sbox_1_and_588 = state_2_41_1_lpi_4 & state_3_41_lpi_3;
  assign Encrypt_Top_sbox_2_and_696 = state_4_4_22_lpi_3 & state_0_22_lpi_6;
  assign Encrypt_Top_sbox_2_and_698 = state_3_22_lpi_3 & state_0_22_lpi_6;
  assign Encrypt_Top_sbox_2_and_700 = state_4_4_40_lpi_3 & state_0_40_lpi_6;
  assign Encrypt_Top_sbox_2_and_702 = state_3_40_lpi_3 & state_0_40_lpi_6;
  assign Encrypt_Top_sbox_1_and_592 = state_2_40_1_lpi_4 & state_3_40_lpi_3;
  assign Encrypt_Top_sbox_2_and_704 = state_4_4_23_lpi_3 & state_0_23_lpi_6;
  assign Encrypt_Top_sbox_2_and_706 = state_3_23_lpi_3 & state_0_23_lpi_6;
  assign Encrypt_Top_sbox_2_and_708 = state_4_4_39_lpi_3 & state_0_39_lpi_6;
  assign Encrypt_Top_sbox_2_and_710 = state_3_39_lpi_3 & state_0_39_lpi_6;
  assign Encrypt_Top_sbox_1_and_596 = state_2_39_1_lpi_4 & state_3_39_lpi_3;
  assign Encrypt_Top_sbox_2_and_716 = state_4_4_38_lpi_3 & state_0_38_lpi_6;
  assign Encrypt_Top_sbox_2_and_718 = state_3_38_lpi_3 & state_0_38_lpi_6;
  assign Encrypt_Top_sbox_1_and_600 = state_2_38_1_lpi_4 & state_3_38_lpi_3;
  assign Encrypt_Top_sbox_2_and_724 = state_4_4_37_lpi_3 & state_0_37_lpi_6;
  assign Encrypt_Top_sbox_2_and_726 = state_3_37_lpi_3 & state_0_37_lpi_6;
  assign Encrypt_Top_sbox_1_and_604 = state_2_37_1_lpi_4 & state_3_37_lpi_3;
  assign Encrypt_Top_sbox_2_and_732 = state_4_4_36_lpi_3 & state_0_36_lpi_6;
  assign Encrypt_Top_sbox_2_and_734 = state_3_36_lpi_3 & state_0_36_lpi_6;
  assign Encrypt_Top_sbox_1_and_608 = state_2_36_1_lpi_4 & state_3_36_lpi_3;
  assign Encrypt_Top_sbox_2_and_740 = state_4_4_35_lpi_3 & state_0_35_lpi_6;
  assign Encrypt_Top_sbox_2_and_742 = state_3_35_lpi_3 & state_0_35_lpi_6;
  assign Encrypt_Top_sbox_1_and_612 = state_2_35_1_lpi_4 & state_3_35_lpi_3;
  assign Encrypt_Top_sbox_2_and_748 = state_4_4_34_lpi_3 & state_0_34_lpi_6;
  assign Encrypt_Top_sbox_2_and_750 = state_3_34_lpi_3 & state_0_34_lpi_6;
  assign Encrypt_Top_sbox_1_and_616 = state_2_34_1_lpi_4 & state_3_34_lpi_3;
  assign Encrypt_Top_sbox_2_and_752 = state_4_4_29_lpi_3 & state_0_29_lpi_6;
  assign Encrypt_Top_sbox_2_and_754 = state_3_29_lpi_3 & state_0_29_lpi_6;
  assign Encrypt_Top_sbox_2_and_756 = state_4_4_33_lpi_3 & state_0_33_lpi_6;
  assign Encrypt_Top_sbox_2_and_758 = state_3_33_lpi_3 & state_0_33_lpi_6;
  assign Encrypt_Top_sbox_1_and_620 = state_2_33_1_lpi_4 & state_3_33_lpi_3;
  assign Encrypt_Top_sbox_2_and_764 = state_4_4_32_lpi_3 & state_0_32_lpi_6;
  assign Encrypt_Top_sbox_2_and_766 = state_3_32_lpi_3 & state_0_32_lpi_6;
  assign Encrypt_Top_sbox_1_and_624 = state_2_32_1_lpi_4 & state_3_32_lpi_3;
  assign Encrypt_Top_sbox_1_and_628 = state_3_0_lpi_3 & state_1_1_31_0_lpi_4_0;
  assign Encrypt_Top_sbox_1_and_630 = state_3_1_lpi_3 & state_1_1_31_0_lpi_4_1;
  assign Encrypt_Top_sbox_1_and_632 = state_3_2_lpi_3 & state_1_1_31_0_lpi_4_2;
  assign Encrypt_Top_sbox_1_and_634 = state_3_3_lpi_3 & state_1_1_31_0_lpi_4_3;
  assign Encrypt_Top_sbox_1_and_636 = state_3_4_lpi_3 & state_1_1_31_0_lpi_4_4;
  assign Encrypt_Top_sbox_1_and_638 = state_3_5_lpi_3 & state_1_1_31_0_lpi_4_5;
  assign Encrypt_Top_sbox_1_and_640 = state_3_6_lpi_3 & state_1_1_31_0_lpi_4_6;
  assign Encrypt_Top_sbox_1_and_642 = state_3_7_lpi_3 & state_1_1_31_0_lpi_4_7;
  assign Encrypt_Top_sbox_1_and_652 = state_3_14_lpi_3 & state_1_1_31_0_lpi_4_14;
  assign Encrypt_Top_sbox_1_and_654 = state_3_15_lpi_3 & state_1_1_31_0_lpi_4_15;
  assign Encrypt_Top_sbox_1_and_656 = state_3_16_lpi_3 & state_1_1_31_0_lpi_4_16;
  assign Encrypt_Top_sbox_1_and_664 = state_3_20_lpi_3 & state_1_1_31_0_lpi_4_20;
  assign Encrypt_Top_sbox_1_and_666 = state_3_21_lpi_3 & state_1_1_31_0_lpi_4_21;
  assign Encrypt_Top_sbox_1_and_694 = state_3_33_lpi_3 & state_1_1_63_32_lpi_4_1;
  assign Encrypt_Top_sbox_1_and_728 = state_3_57_lpi_3 & state_1_1_63_32_lpi_4_25;
  assign Encrypt_Top_sbox_1_and_734 = state_3_60_lpi_3 & state_1_1_63_32_lpi_4_28;
  assign Encrypt_Top_sbox_1_and_756 = state_4_4_0_lpi_3 & state_3_0_lpi_3;
  assign Encrypt_Top_sbox_1_and_758 = state_4_4_1_lpi_3 & state_3_1_lpi_3;
  assign Encrypt_Top_sbox_1_and_760 = state_4_4_2_lpi_3 & state_3_2_lpi_3;
  assign Encrypt_Top_sbox_1_and_762 = state_4_4_3_lpi_3 & state_3_3_lpi_3;
  assign Encrypt_Top_sbox_1_and_764 = state_4_4_4_lpi_3 & state_3_4_lpi_3;
  assign Encrypt_Top_sbox_1_and_766 = state_4_4_5_lpi_3 & state_3_5_lpi_3;
  assign Encrypt_Top_sbox_1_and_768 = state_4_4_6_lpi_3 & state_3_6_lpi_3;
  assign Encrypt_Top_sbox_1_and_770 = state_4_4_7_lpi_3 & state_3_7_lpi_3;
  assign Encrypt_Top_sbox_1_and_784 = state_4_4_16_lpi_3 & state_3_16_lpi_3;
  assign Encrypt_Top_sbox_1_and_786 = state_4_4_17_lpi_3 & state_3_17_lpi_3;
  assign Encrypt_Top_sbox_1_and_788 = state_4_4_18_lpi_3 & state_3_18_lpi_3;
  assign Encrypt_Top_sbox_1_and_790 = state_4_4_19_lpi_3 & state_3_19_lpi_3;
  assign Encrypt_Top_sbox_1_and_792 = state_4_4_20_lpi_3 & state_3_20_lpi_3;
  assign Encrypt_Top_sbox_1_and_796 = state_4_4_22_lpi_3 & state_3_22_lpi_3;
  assign Encrypt_Top_sbox_1_and_798 = state_4_4_23_lpi_3 & state_3_23_lpi_3;
  assign Encrypt_Top_sbox_1_and_800 = state_4_4_24_lpi_3 & state_3_24_lpi_3;
  assign Encrypt_Top_sbox_1_and_802 = state_4_4_25_lpi_3 & state_3_25_lpi_3;
  assign Encrypt_Top_sbox_1_and_808 = state_4_4_28_lpi_3 & state_3_28_lpi_3;
  assign Encrypt_Top_sbox_1_and_816 = state_4_4_32_lpi_3 & state_3_32_lpi_3;
  assign Encrypt_Top_sbox_1_and_818 = state_4_4_33_lpi_3 & state_3_33_lpi_3;
  assign Encrypt_Top_sbox_1_and_820 = state_4_4_34_lpi_3 & state_3_34_lpi_3;
  assign Encrypt_Top_sbox_1_and_822 = state_4_4_35_lpi_3 & state_3_35_lpi_3;
  assign Encrypt_Top_sbox_1_and_824 = state_4_4_36_lpi_3 & state_3_36_lpi_3;
  assign Encrypt_Top_sbox_1_and_826 = state_4_4_37_lpi_3 & state_3_37_lpi_3;
  assign Encrypt_Top_sbox_1_and_828 = state_4_4_38_lpi_3 & state_3_38_lpi_3;
  assign Encrypt_Top_sbox_1_and_830 = state_4_4_39_lpi_3 & state_3_39_lpi_3;
  assign Encrypt_Top_sbox_1_and_832 = state_4_4_40_lpi_3 & state_3_40_lpi_3;
  assign Encrypt_Top_sbox_1_and_834 = state_4_4_41_lpi_3 & state_3_41_lpi_3;
  assign Encrypt_Top_sbox_1_and_836 = state_4_4_42_lpi_3 & state_3_42_lpi_3;
  assign Encrypt_Top_sbox_1_and_838 = state_4_4_43_lpi_3 & state_3_43_lpi_3;
  assign Encrypt_Top_sbox_1_and_840 = state_4_4_44_lpi_3 & state_3_44_lpi_3;
  assign Encrypt_Top_sbox_1_and_842 = state_4_4_45_lpi_3 & state_3_45_lpi_3;
  assign Encrypt_Top_sbox_1_and_844 = state_4_4_46_lpi_3 & state_3_46_lpi_3;
  assign Encrypt_Top_sbox_1_and_846 = state_4_4_47_lpi_3 & state_3_47_lpi_3;
  assign Encrypt_Top_sbox_1_and_848 = state_4_4_48_lpi_3 & state_3_48_lpi_3;
  assign Encrypt_Top_sbox_1_and_850 = state_4_4_49_lpi_3 & state_3_49_lpi_3;
  assign Encrypt_Top_sbox_1_and_852 = state_4_4_50_lpi_3 & state_3_50_lpi_3;
  assign Encrypt_Top_sbox_1_and_854 = state_4_4_51_lpi_3 & state_3_51_lpi_3;
  assign Encrypt_Top_sbox_1_and_856 = state_4_4_52_lpi_3 & state_3_52_lpi_3;
  assign Encrypt_Top_sbox_1_and_858 = state_4_4_53_lpi_3 & state_3_53_lpi_3;
  assign Encrypt_Top_sbox_1_and_860 = state_4_4_54_lpi_3 & state_3_54_lpi_3;
  assign Encrypt_Top_sbox_1_and_862 = state_4_4_55_lpi_3 & state_3_55_lpi_3;
  assign Encrypt_Top_sbox_1_and_864 = state_4_4_56_lpi_3 & state_3_56_lpi_3;
  assign Encrypt_Top_sbox_1_and_866 = state_4_4_57_lpi_3 & state_3_57_lpi_3;
  assign Encrypt_Top_sbox_1_and_868 = state_4_4_58_lpi_3 & state_3_58_lpi_3;
  assign Encrypt_Top_sbox_1_and_870 = state_4_4_59_lpi_3 & state_3_59_lpi_3;
  assign Encrypt_Top_sbox_1_and_872 = state_4_4_60_lpi_3 & state_3_60_lpi_3;
  assign Encrypt_Top_sbox_1_and_874 = state_4_4_61_lpi_3 & state_3_61_lpi_3;
  assign Encrypt_Top_sbox_1_and_876 = state_4_4_62_lpi_3 & state_3_62_lpi_3;
  assign Encrypt_Top_sbox_1_and_878 = state_4_4_63_lpi_3 & state_3_63_lpi_3;
  assign Encrypt_Top_sbox_1_and_880 = state_4_4_8_lpi_3 & state_3_8_lpi_3;
  assign Encrypt_Top_sbox_1_and_882 = state_4_4_9_lpi_3 & state_3_9_lpi_3;
  assign operator_33_true_1_operator_33_true_1_and_tmp = (({ADLEN_i_7_0_sva_6_4 ,
      ADLEN_i_7_0_sva_3_0}) == (z_out[6:0])) & (z_out[8:7]==2'b00);
  assign or_dcpl_9 = (z_out_2[7]) | operator_33_true_1_operator_33_true_1_and_tmp;
  assign and_24_cse = (fsm_output[11]) | (fsm_output[4]);
  assign and_90_cse = (~ z_out_1_2) & (fsm_output[11]);
  assign and_94_cse = (~ z_out_1_2) & (fsm_output[14]);
  assign and_738_cse = (~((z_out_2[7]) | operator_33_true_1_operator_33_true_1_and_tmp))
      & (fsm_output[13]);
  assign and_740_cse = (~ z_out_1_2) & (fsm_output[1]);
  assign or_tmp_382 = and_24_cse | and_39_cse;
  assign and_885_cse = or_dcpl_9 & (fsm_output[13]);
  assign or_tmp_913 = and_21_cse | (fsm_output[4]);
  assign or_tmp_1693 = and_24_cse | (fsm_output[14]);
  assign ADLEN_i_7_0_sva_6_0_mx0c3 = and_885_cse | (z_out_1_2 & (fsm_output[1]))
      | (fsm_output[0]) | (fsm_output[14]);
  assign xor_cse_1 = state_1_1_63_32_lpi_4_19 ^ (state_4_4_51_lpi_3 & state_1_1_63_32_lpi_4_19)
      ^ state_3_51_lpi_3 ^ (state_1_1_63_32_lpi_4_19 & state_0_51_lpi_6);
  assign xor_cse = state_0_51_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_51_sva_1 ^ xor_cse_1
      ^ state_2_51_1_lpi_4;
  assign xor_cse_3 = state_2_60_1_lpi_4 ^ state_0_60_lpi_6 ^ state_3_60_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_60_sva_1;
  assign xor_cse_4 = state_1_1_63_32_lpi_4_0 ^ (state_4_4_32_lpi_3 & state_1_1_63_32_lpi_4_0)
      ^ state_3_32_lpi_3 ^ (state_1_1_63_32_lpi_4_0 & state_0_32_lpi_6);
  assign xor_cse_5 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_2_and_2_cse_60_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_32_sva_1;
  assign ciphertext_32_sva_mx0w2 = xor_cse ^ xor_cse_3 ^ xor_cse_4 ^ xor_cse_5 ^
      plaintext_63_32_sva_0 ^ state_2_32_1_lpi_4 ^ state_0_32_lpi_6;
  assign xor_cse_8 = state_2_42_1_lpi_4 ^ state_0_42_lpi_6 ^ state_3_42_lpi_3 ^ state_4_4_42_lpi_3;
  assign xor_cse_7 = xor_cse_8 ^ Encrypt_Top_sbox_2_and_684 ^ Encrypt_Top_sbox_2_and_686
      ^ Encrypt_Top_sbox_2_and_766;
  assign xor_cse_10 = state_2_49_1_lpi_4 ^ state_0_49_lpi_6 ^ state_3_49_lpi_3 ^
      state_4_4_49_lpi_3;
  assign xor_cse_11 = state_2_32_1_lpi_4 ^ state_0_32_lpi_6 ^ state_3_32_lpi_3 ^
      state_4_4_32_lpi_3;
  assign xor_cse_12 = Encrypt_Top_sbox_2_and_628 ^ Encrypt_Top_sbox_2_and_630 ^ state_1_1_63_32_lpi_4_22
      ^ Encrypt_Top_sbox_2_and_764;
  assign xor_cse_15 = state_1_1_63_32_lpi_4_20 ^ (state_4_4_52_lpi_3 & state_1_1_63_32_lpi_4_20)
      ^ state_3_52_lpi_3 ^ (state_1_1_63_32_lpi_4_20 & state_0_52_lpi_6);
  assign xor_cse_14 = state_0_52_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_52_sva_1 ^
      xor_cse_15 ^ state_2_52_1_lpi_4;
  assign xor_cse_17 = state_2_61_1_lpi_4 ^ state_0_61_lpi_6 ^ state_3_61_lpi_3 ^
      Encrypt_Top_sbox_1_and_cse_61_sva_1;
  assign xor_cse_18 = state_1_1_63_32_lpi_4_1 ^ (state_4_4_33_lpi_3 & state_1_1_63_32_lpi_4_1)
      ^ state_3_33_lpi_3 ^ (state_1_1_63_32_lpi_4_1 & state_0_33_lpi_6);
  assign xor_cse_19 = state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_1_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_61_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1;
  assign ciphertext_33_sva_mx0w2 = xor_cse_14 ^ xor_cse_17 ^ xor_cse_18 ^ xor_cse_19
      ^ plaintext_63_32_sva_1 ^ state_2_33_1_lpi_4 ^ state_0_33_lpi_6;
  assign xor_cse_22 = state_2_43_1_lpi_4 ^ state_0_43_lpi_6 ^ state_3_43_lpi_3 ^
      state_4_4_43_lpi_3;
  assign xor_cse_21 = xor_cse_22 ^ Encrypt_Top_sbox_2_and_676 ^ Encrypt_Top_sbox_2_and_678
      ^ Encrypt_Top_sbox_2_and_758;
  assign xor_cse_24 = state_2_50_1_lpi_4 ^ state_0_50_lpi_6 ^ state_3_50_lpi_3 ^
      state_4_4_50_lpi_3;
  assign xor_cse_25 = state_2_33_1_lpi_4 ^ state_0_33_lpi_6 ^ state_3_33_lpi_3 ^
      state_4_4_33_lpi_3;
  assign xor_cse_26 = state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_2_and_620 ^ Encrypt_Top_sbox_2_and_622
      ^ Encrypt_Top_sbox_2_and_756;
  assign xor_cse_28 = state_2_62_1_lpi_4 ^ state_0_62_lpi_6 ^ state_3_62_lpi_3 ^
      Encrypt_Top_sbox_1_and_cse_62_sva_1;
  assign xor_cse_29 = state_1_1_63_32_lpi_4_21 ^ (state_4_4_53_lpi_3 & state_1_1_63_32_lpi_4_21)
      ^ state_3_53_lpi_3 ^ (state_1_1_63_32_lpi_4_21 & state_0_53_lpi_6);
  assign xor_cse_30 = state_1_1_63_32_lpi_4_2 ^ (state_4_4_34_lpi_3 & state_1_1_63_32_lpi_4_2)
      ^ state_3_34_lpi_3 ^ (state_1_1_63_32_lpi_4_2 & state_0_34_lpi_6);
  assign xor_cse_31 = state_1_1_63_32_lpi_4_30 ^ Encrypt_Top_sbox_1_and_1_cse_62_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_62_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1;
  assign xor_cse_32 = state_2_34_1_lpi_4 ^ state_0_34_lpi_6 ^ state_2_53_1_lpi_4
      ^ state_0_53_lpi_6;
  assign ciphertext_34_sva_mx0w2 = xor_cse_28 ^ xor_cse_29 ^ xor_cse_30 ^ xor_cse_31
      ^ xor_cse_32 ^ plaintext_63_32_sva_2 ^ Encrypt_Top_sbox_1_and_1_cse_53_sva_1;
  assign xor_cse_35 = state_2_44_1_lpi_4 ^ state_0_44_lpi_6 ^ state_3_44_lpi_3 ^
      state_4_4_44_lpi_3;
  assign xor_cse_34 = xor_cse_35 ^ Encrypt_Top_sbox_2_and_668 ^ Encrypt_Top_sbox_2_and_670
      ^ state_1_1_63_32_lpi_4_18;
  assign xor_cse_37 = state_2_51_1_lpi_4 ^ state_0_51_lpi_6 ^ state_3_51_lpi_3 ^
      state_4_4_51_lpi_3;
  assign xor_cse_38 = state_2_34_1_lpi_4 ^ state_0_34_lpi_6 ^ state_3_34_lpi_3 ^
      state_4_4_34_lpi_3;
  assign xor_cse_39 = state_1_1_63_32_lpi_4_24 ^ Encrypt_Top_sbox_2_and_612 ^ Encrypt_Top_sbox_2_and_614
      ^ Encrypt_Top_sbox_2_and_748;
  assign xor_cse_42 = state_1_1_63_32_lpi_4_31 ^ (state_4_4_63_lpi_3 & state_1_1_63_32_lpi_4_31)
      ^ state_3_63_lpi_3 ^ (state_1_1_63_32_lpi_4_31 & state_0_63_lpi_6);
  assign xor_cse_41 = state_0_63_lpi_6 ^ state_2_63_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_63_sva_1
      ^ xor_cse_42;
  assign xor_cse_44 = state_1_1_63_32_lpi_4_22 ^ (state_4_4_54_lpi_3 & state_1_1_63_32_lpi_4_22)
      ^ state_3_54_lpi_3 ^ (state_1_1_63_32_lpi_4_22 & state_0_54_lpi_6);
  assign xor_cse_43 = state_2_54_1_lpi_4 ^ state_0_54_lpi_6 ^ xor_cse_44;
  assign xor_cse_46 = state_1_1_63_32_lpi_4_3 ^ (state_4_4_35_lpi_3 & state_1_1_63_32_lpi_4_3)
      ^ state_3_35_lpi_3 ^ (state_1_1_63_32_lpi_4_3 & state_0_35_lpi_6);
  assign xor_cse_47 = state_2_35_1_lpi_4 ^ state_0_35_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_35_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1;
  assign ciphertext_35_sva_mx0w2 = xor_cse_41 ^ xor_cse_43 ^ plaintext_63_32_sva_3
      ^ xor_cse_46 ^ xor_cse_47;
  assign xor_cse_49 = state_2_45_1_lpi_4 ^ state_0_45_lpi_6 ^ state_3_45_lpi_3 ^
      state_4_4_45_lpi_3;
  assign xor_cse_48 = xor_cse_49 ^ Encrypt_Top_sbox_2_and_662 ^ Encrypt_Top_sbox_2_and_660
      ^ Encrypt_Top_sbox_2_and_742;
  assign xor_cse_51 = state_2_52_1_lpi_4 ^ state_0_52_lpi_6 ^ state_3_52_lpi_3 ^
      state_4_4_52_lpi_3;
  assign xor_cse_52 = state_2_35_1_lpi_4 ^ state_0_35_lpi_6 ^ state_3_35_lpi_3 ^
      state_4_4_35_lpi_3;
  assign xor_cse_53 = state_1_1_63_32_lpi_4_25 ^ Encrypt_Top_sbox_2_and_604 ^ Encrypt_Top_sbox_2_and_606
      ^ Encrypt_Top_sbox_2_and_740;
  assign xor_cse_56 = state_1_1_31_0_lpi_4_0 ^ (state_4_4_0_lpi_3 & state_1_1_31_0_lpi_4_0)
      ^ state_3_0_lpi_3 ^ (state_1_1_31_0_lpi_4_0 & state_0_0_lpi_6);
  assign xor_cse_57 = state_1_1_63_32_lpi_4_23 ^ (state_4_4_55_lpi_3 & state_1_1_63_32_lpi_4_23)
      ^ state_3_55_lpi_3 ^ (state_1_1_63_32_lpi_4_23 & state_0_55_lpi_6);
  assign xor_cse_55 = xor_cse_56 ^ state_0_36_lpi_6 ^ state_2_36_1_lpi_4 ^ xor_cse_57;
  assign xor_cse_59 = state_1_1_63_32_lpi_4_4 ^ (state_4_4_36_lpi_3 & state_1_1_63_32_lpi_4_4)
      ^ state_3_36_lpi_3 ^ (state_1_1_63_32_lpi_4_4 & state_0_36_lpi_6);
  assign xor_cse_60 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]) ^ state_0_0_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_0_sva_1 ^ state_2_0_1_lpi_6;
  assign xor_cse_61 = state_2_55_1_lpi_4 ^ state_0_55_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_55_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_36_sva_1;
  assign ciphertext_36_sva_mx0w2 = xor_cse_55 ^ plaintext_63_32_sva_4 ^ xor_cse_59
      ^ xor_cse_60 ^ xor_cse_61;
  assign xor_cse_63 = state_2_46_1_lpi_4 ^ state_0_46_lpi_6 ^ state_3_46_lpi_3 ^
      state_4_4_46_lpi_3;
  assign xor_cse_62 = xor_cse_63 ^ Encrypt_Top_sbox_2_and_654 ^ Encrypt_Top_sbox_2_and_652
      ^ Encrypt_Top_sbox_2_and_734;
  assign xor_cse_65 = state_2_53_1_lpi_4 ^ state_0_53_lpi_6 ^ state_3_53_lpi_3 ^
      state_4_4_53_lpi_3;
  assign xor_cse_66 = state_2_36_1_lpi_4 ^ state_0_36_lpi_6 ^ state_3_36_lpi_3 ^
      state_4_4_36_lpi_3;
  assign xor_cse_67 = state_1_1_63_32_lpi_4_26 ^ Encrypt_Top_sbox_2_and_596 ^ Encrypt_Top_sbox_2_and_598
      ^ Encrypt_Top_sbox_2_and_732;
  assign xor_cse_70 = state_1_1_31_0_lpi_4_1 ^ (state_4_4_1_lpi_3 & state_1_1_31_0_lpi_4_1)
      ^ state_3_1_lpi_3 ^ (state_1_1_31_0_lpi_4_1 & state_0_1_lpi_6);
  assign xor_cse_71 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]) ^ state_0_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_1_sva_1 ^ state_2_1_1_lpi_6;
  assign xor_cse_69 = xor_cse_70 ^ xor_cse_71 ^ state_2_37_1_lpi_4 ^ state_0_37_lpi_6;
  assign xor_cse_73 = state_1_1_63_32_lpi_4_24 ^ (state_4_4_56_lpi_3 & state_1_1_63_32_lpi_4_24)
      ^ state_3_56_lpi_3 ^ (state_1_1_63_32_lpi_4_24 & state_0_56_lpi_6);
  assign xor_cse_74 = state_1_1_63_32_lpi_4_5 ^ (state_4_4_37_lpi_3 & state_1_1_63_32_lpi_4_5)
      ^ state_3_37_lpi_3 ^ (state_1_1_63_32_lpi_4_5 & state_0_37_lpi_6);
  assign xor_cse_75 = state_2_56_1_lpi_4 ^ state_0_56_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_56_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1;
  assign ciphertext_37_sva_mx0w2 = xor_cse_69 ^ plaintext_63_32_sva_5 ^ xor_cse_73
      ^ xor_cse_74 ^ xor_cse_75;
  assign xor_cse_77 = state_2_47_1_lpi_4 ^ state_0_47_lpi_6 ^ state_3_47_lpi_3 ^
      state_4_4_47_lpi_3;
  assign xor_cse_76 = xor_cse_77 ^ Encrypt_Top_sbox_2_and_646 ^ Encrypt_Top_sbox_2_and_644
      ^ Encrypt_Top_sbox_2_and_726;
  assign xor_cse_79 = state_2_54_1_lpi_4 ^ state_0_54_lpi_6 ^ state_3_54_lpi_3 ^
      state_4_4_54_lpi_3;
  assign xor_cse_80 = state_2_37_1_lpi_4 ^ state_0_37_lpi_6 ^ state_3_37_lpi_3 ^
      state_4_4_37_lpi_3;
  assign xor_cse_81 = state_1_1_63_32_lpi_4_27 ^ Encrypt_Top_sbox_2_and_588 ^ Encrypt_Top_sbox_2_and_590
      ^ Encrypt_Top_sbox_2_and_724;
  assign xor_cse_84 = state_1_1_31_0_lpi_4_2 ^ (state_4_4_2_lpi_3 & state_1_1_31_0_lpi_4_2)
      ^ state_3_2_lpi_3 ^ (state_1_1_31_0_lpi_4_2 & state_0_2_lpi_6);
  assign xor_cse_85 = state_1_1_63_32_lpi_4_25 ^ (state_4_4_57_lpi_3 & state_1_1_63_32_lpi_4_25)
      ^ state_3_57_lpi_3 ^ (state_1_1_63_32_lpi_4_25 & state_0_57_lpi_6);
  assign xor_cse_83 = xor_cse_84 ^ state_2_38_1_lpi_4 ^ state_0_38_lpi_6 ^ xor_cse_85;
  assign xor_cse_87 = state_1_1_63_32_lpi_4_6 ^ (state_4_4_38_lpi_3 & state_1_1_63_32_lpi_4_6)
      ^ state_3_38_lpi_3 ^ (state_1_1_63_32_lpi_4_6 & state_0_38_lpi_6);
  assign xor_cse_88 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]) ^ state_0_2_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_2_sva_1 ^ state_2_2_1_lpi_6;
  assign xor_cse_89 = state_2_57_1_lpi_4 ^ state_0_57_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1;
  assign ciphertext_38_sva_mx0w2 = xor_cse_83 ^ plaintext_63_32_sva_6 ^ xor_cse_87
      ^ xor_cse_88 ^ xor_cse_89;
  assign xor_cse_91 = state_2_55_1_lpi_4 ^ state_0_55_lpi_6 ^ state_3_55_lpi_3 ^
      state_4_4_55_lpi_3;
  assign xor_cse_92 = state_2_38_1_lpi_4 ^ state_0_38_lpi_6 ^ state_3_38_lpi_3 ^
      state_4_4_38_lpi_3;
  assign xor_cse_90 = xor_cse_91 ^ Encrypt_Top_sbox_2_and_718 ^ xor_cse_92 ^ state_1_1_63_32_lpi_4_12;
  assign xor_cse_94 = state_2_48_1_lpi_4 ^ state_0_48_lpi_6 ^ state_3_48_lpi_3 ^
      state_4_4_48_lpi_3;
  assign xor_cse_95 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_2_and_580 ^ Encrypt_Top_sbox_2_and_582
      ^ Encrypt_Top_sbox_2_and_716;
  assign xor_cse_98 = state_1_1_63_32_lpi_4_7 ^ (state_4_4_39_lpi_3 & state_1_1_63_32_lpi_4_7)
      ^ state_3_39_lpi_3 ^ (state_1_1_63_32_lpi_4_7 & state_0_39_lpi_6);
  assign xor_cse_97 = state_2_39_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_39_sva_1
      ^ xor_cse_98 ^ Encrypt_Top_sbox_1_and_1_cse_58_sva_1;
  assign xor_cse_100 = state_1_1_63_32_lpi_4_26 ^ (state_4_4_58_lpi_3 & state_1_1_63_32_lpi_4_26)
      ^ state_3_58_lpi_3 ^ (state_1_1_63_32_lpi_4_26 & state_0_58_lpi_6);
  assign xor_cse_99 = state_0_58_lpi_6 ^ xor_cse_100 ^ state_2_58_1_lpi_4 ^ state_0_39_lpi_6;
  assign xor_cse_102 = state_1_1_31_0_lpi_4_3 ^ (state_4_4_3_lpi_3 & state_1_1_31_0_lpi_4_3)
      ^ state_3_3_lpi_3 ^ (state_1_1_31_0_lpi_4_3 & state_0_3_lpi_6);
  assign xor_cse_103 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]) ^ state_0_3_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_3_sva_1 ^ state_2_3_1_lpi_6;
  assign ciphertext_39_sva_mx0w2 = xor_cse_97 ^ xor_cse_99 ^ plaintext_63_32_sva_7
      ^ xor_cse_102 ^ xor_cse_103;
  assign xor_cse_104 = xor_cse_10 ^ Encrypt_Top_sbox_2_and_628 ^ Encrypt_Top_sbox_2_and_630
      ^ Encrypt_Top_sbox_2_and_710;
  assign xor_cse_106 = state_2_56_1_lpi_4 ^ state_0_56_lpi_6 ^ state_3_56_lpi_3 ^
      state_4_4_56_lpi_3;
  assign xor_cse_107 = state_2_39_1_lpi_4 ^ state_0_39_lpi_6 ^ state_3_39_lpi_3 ^
      state_4_4_39_lpi_3;
  assign xor_cse_108 = state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_2_and_572 ^ Encrypt_Top_sbox_2_and_574
      ^ Encrypt_Top_sbox_2_and_708;
  assign xor_cse_111 = state_1_1_31_0_lpi_4_4 ^ (state_4_4_4_lpi_3 & state_1_1_31_0_lpi_4_4)
      ^ state_3_4_lpi_3 ^ (state_1_1_31_0_lpi_4_4 & state_0_4_lpi_6);
  assign xor_cse_110 = xor_cse_111 ^ state_0_59_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_40_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_59_sva_1;
  assign xor_cse_113 = state_1_1_63_32_lpi_4_8 ^ (state_4_4_40_lpi_3 & state_1_1_63_32_lpi_4_8)
      ^ state_3_40_lpi_3 ^ (state_1_1_63_32_lpi_4_8 & state_0_40_lpi_6);
  assign xor_cse_112 = state_2_40_1_lpi_4 ^ state_0_40_lpi_6 ^ xor_cse_113 ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1;
  assign xor_cse_115 = state_1_1_63_32_lpi_4_27 ^ state_2_59_1_lpi_4 ^ Encrypt_Top_sbox_1_and_cse_59_sva_1
      ^ state_3_59_lpi_3;
  assign xor_cse_116 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]) ^ state_0_4_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_4_sva_1 ^ state_2_4_1_lpi_6;
  assign ciphertext_40_sva_mx0w2 = xor_cse_110 ^ xor_cse_112 ^ plaintext_63_32_sva_8
      ^ xor_cse_115 ^ xor_cse_116;
  assign xor_cse_117 = xor_cse_24 ^ Encrypt_Top_sbox_2_and_622 ^ Encrypt_Top_sbox_2_and_620
      ^ Encrypt_Top_sbox_2_and_702;
  assign xor_cse_119 = state_2_57_1_lpi_4 ^ state_0_57_lpi_6 ^ state_3_57_lpi_3 ^
      state_4_4_57_lpi_3;
  assign xor_cse_120 = state_2_40_1_lpi_4 ^ state_0_40_lpi_6 ^ state_3_40_lpi_3 ^
      state_4_4_40_lpi_3;
  assign xor_cse_121 = state_1_1_63_32_lpi_4_3 ^ Encrypt_Top_sbox_2_and_566 ^ Encrypt_Top_sbox_2_and_564
      ^ Encrypt_Top_sbox_2_and_700;
  assign xor_cse_124 = state_1_1_31_0_lpi_4_5 ^ (state_4_4_5_lpi_3 & state_1_1_31_0_lpi_4_5)
      ^ state_3_5_lpi_3 ^ (state_1_1_31_0_lpi_4_5 & state_0_5_lpi_6);
  assign xor_cse_125 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]) ^ state_2_5_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_5_sva_1 ^ state_0_5_lpi_6;
  assign xor_cse_123 = xor_cse_124 ^ xor_cse_125 ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1
      ^ state_0_41_lpi_6;
  assign xor_cse_127 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_2_and_2_cse_60_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1 ^ Encrypt_Top_sbox_1_and_cse_41_sva_1;
  assign xor_cse_128 = state_1_1_63_32_lpi_4_9 ^ Encrypt_Top_sbox_1_and_1_cse_41_sva_1
      ^ state_3_41_lpi_3 ^ state_2_41_1_lpi_4;
  assign ciphertext_41_sva_mx0w2 = xor_cse_123 ^ plaintext_63_32_sva_9 ^ xor_cse_3
      ^ xor_cse_127 ^ xor_cse_128;
  assign xor_cse_130 = state_2_41_1_lpi_4 ^ state_0_41_lpi_6 ^ state_3_41_lpi_3 ^
      state_4_4_41_lpi_3;
  assign xor_cse_129 = xor_cse_130 ^ Encrypt_Top_sbox_2_and_694 ^ Encrypt_Top_sbox_2_and_612
      ^ Encrypt_Top_sbox_2_and_614;
  assign xor_cse_132 = state_2_58_1_lpi_4 ^ state_0_58_lpi_6 ^ state_3_58_lpi_3 ^
      state_4_4_58_lpi_3;
  assign xor_cse_133 = state_1_1_63_32_lpi_4_30 ^ Encrypt_Top_sbox_2_and_558 ^ Encrypt_Top_sbox_2_and_556
      ^ Encrypt_Top_sbox_2_and_692;
  assign xor_cse_136 = state_1_1_31_0_lpi_4_6 ^ (state_4_4_6_lpi_3 & state_1_1_31_0_lpi_4_6)
      ^ state_3_6_lpi_3 ^ (state_1_1_31_0_lpi_4_6 & state_0_6_lpi_6);
  assign xor_cse_137 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]) ^ state_2_6_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_6_sva_1 ^ state_0_6_lpi_6;
  assign xor_cse_135 = xor_cse_136 ^ xor_cse_137 ^ Encrypt_Top_sbox_2_and_2_cse_42_sva_1
      ^ state_0_42_lpi_6;
  assign xor_cse_139 = state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_1_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_61_sva_1 ^ Encrypt_Top_sbox_1_and_cse_42_sva_1;
  assign xor_cse_140 = state_1_1_63_32_lpi_4_10 ^ state_2_42_1_lpi_4 ^ state_3_42_lpi_3
      ^ Encrypt_Top_sbox_1_and_1_cse_42_sva_1;
  assign ciphertext_42_sva_mx0w2 = xor_cse_135 ^ plaintext_63_32_sva_10 ^ xor_cse_17
      ^ xor_cse_139 ^ xor_cse_140;
  assign xor_cse_142 = state_2_59_1_lpi_4 ^ state_0_59_lpi_6 ^ state_3_59_lpi_3 ^
      state_4_4_59_lpi_3;
  assign xor_cse_141 = xor_cse_142 ^ Encrypt_Top_sbox_2_and_550 ^ state_1_1_63_32_lpi_4_31
      ^ Encrypt_Top_sbox_2_and_548;
  assign xor_cse_143 = xor_cse_51 ^ Encrypt_Top_sbox_2_and_606 ^ xor_cse_8;
  assign xor_cse_145 = state_1_1_63_32_lpi_4_16 ^ Encrypt_Top_sbox_2_and_684 ^ Encrypt_Top_sbox_2_and_686
      ^ Encrypt_Top_sbox_2_and_604;
  assign xor_cse_148 = state_1_1_31_0_lpi_4_7 ^ (state_4_4_7_lpi_3 & state_1_1_31_0_lpi_4_7)
      ^ state_3_7_lpi_3 ^ (state_1_1_31_0_lpi_4_7 & state_0_7_lpi_6);
  assign xor_cse_149 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]) ^ state_2_7_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_7_sva_1 ^ state_0_7_lpi_6;
  assign xor_cse_147 = xor_cse_148 ^ xor_cse_149 ^ state_2_43_1_lpi_4 ^ state_0_43_lpi_6;
  assign xor_cse_151 = state_1_1_63_32_lpi_4_11 ^ (state_4_4_43_lpi_3 & state_1_1_63_32_lpi_4_11)
      ^ state_3_43_lpi_3 ^ (state_1_1_63_32_lpi_4_11 & state_0_43_lpi_6);
  assign xor_cse_152 = state_1_1_63_32_lpi_4_30 ^ Encrypt_Top_sbox_1_and_1_cse_62_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_62_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_43_sva_1;
  assign ciphertext_43_sva_mx0w2 = xor_cse_147 ^ plaintext_63_32_sva_11 ^ xor_cse_28
      ^ xor_cse_151 ^ xor_cse_152;
  assign xor_cse_154 = state_2_60_1_lpi_4 ^ state_0_60_lpi_6 ^ state_3_60_lpi_3 ^
      state_4_4_60_lpi_3;
  assign xor_cse_153 = xor_cse_154 ^ Encrypt_Top_sbox_2_and_542 ^ state_1_1_63_32_lpi_4_4
      ^ Encrypt_Top_sbox_2_and_540;
  assign xor_cse_156 = state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_2_and_676 ^ Encrypt_Top_sbox_2_and_678
      ^ Encrypt_Top_sbox_2_and_596;
  assign xor_cse_159 = state_1_1_31_0_lpi_4_8 ^ (state_4_4_8_lpi_3 & state_1_1_31_0_lpi_4_8)
      ^ state_3_8_lpi_3 ^ (state_1_1_31_0_lpi_4_8 & state_0_8_lpi_6);
  assign xor_cse_160 = state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_1_and_1_cse_44_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_44_sva_1 ^ state_3_44_lpi_3;
  assign xor_cse_161 = state_2_8_1_lpi_4 ^ state_0_8_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_8_sva_1
      ^ state_2_44_1_lpi_4;
  assign ciphertext_44_sva_mx0w2 = xor_cse_41 ^ xor_cse_159 ^ xor_cse_160 ^ xor_cse_161
      ^ plaintext_63_32_sva_12 ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1 ^ state_0_44_lpi_6;
  assign xor_cse_164 = state_2_61_1_lpi_4 ^ state_0_61_lpi_6 ^ state_3_61_lpi_3 ^
      state_4_4_61_lpi_3;
  assign xor_cse_163 = xor_cse_164 ^ Encrypt_Top_sbox_2_and_534 ^ Encrypt_Top_sbox_2_and_588
      ^ Encrypt_Top_sbox_2_and_590;
  assign xor_cse_168 = state_1_1_63_32_lpi_4_13 ^ (state_4_4_45_lpi_3 & state_1_1_63_32_lpi_4_13)
      ^ state_3_45_lpi_3 ^ (state_1_1_63_32_lpi_4_13 & state_0_45_lpi_6);
  assign xor_cse_167 = state_2_45_1_lpi_4 ^ state_0_45_lpi_6 ^ xor_cse_168 ^ xor_cse_56;
  assign xor_cse_170 = state_1_1_31_0_lpi_4_9 ^ (state_4_4_9_lpi_3 & state_1_1_31_0_lpi_4_9)
      ^ state_3_9_lpi_3 ^ (state_1_1_31_0_lpi_4_9 & state_0_9_lpi_6);
  assign xor_cse_171 = state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_9_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_45_sva_1;
  assign ciphertext_45_sva_mx0w2 = xor_cse_167 ^ plaintext_63_32_sva_13 ^ xor_cse_170
      ^ xor_cse_60 ^ xor_cse_171;
  assign xor_cse_172 = state_1_1_63_32_lpi_4_28 ^ xor_cse_91 ^ Encrypt_Top_sbox_2_and_580
      ^ Encrypt_Top_sbox_2_and_582;
  assign xor_cse_174 = state_2_62_1_lpi_4 ^ state_0_62_lpi_6 ^ state_3_62_lpi_3 ^
      state_4_4_62_lpi_3;
  assign xor_cse_175 = state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_2_and_524 ^ Encrypt_Top_sbox_2_and_526
      ^ Encrypt_Top_sbox_2_and_660;
  assign xor_cse_178 = state_2_10_1_lpi_4 ^ state_0_10_lpi_6 ^ state_3_10_lpi_3 ^
      state_1_1_31_0_lpi_4_10;
  assign xor_cse_177 = xor_cse_178 ^ state_0_46_lpi_6 ^ xor_cse_70 ^ Encrypt_Top_sbox_1_and_cse_10_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_10_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_10_sva_1
      ^ state_2_46_1_lpi_4;
  assign xor_cse_181 = state_1_1_63_32_lpi_4_14 ^ (state_4_4_46_lpi_3 & state_1_1_63_32_lpi_4_14)
      ^ state_3_46_lpi_3 ^ (state_1_1_63_32_lpi_4_14 & state_0_46_lpi_6);
  assign ciphertext_46_sva_mx0w2 = xor_cse_177 ^ xor_cse_181 ^ xor_cse_71 ^ plaintext_63_32_sva_14
      ^ Encrypt_Top_sbox_1_and_1_cse_46_sva_1;
  assign xor_cse_183 = xor_cse_106 ^ Encrypt_Top_sbox_2_and_574 ^ Encrypt_Top_sbox_2_and_572
      ^ state_1_1_63_32_lpi_4_29;
  assign xor_cse_185 = state_2_63_1_lpi_4 ^ state_0_63_lpi_6 ^ state_3_63_lpi_3 ^
      state_4_4_63_lpi_3;
  assign xor_cse_186 = state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_2_and_518 ^ Encrypt_Top_sbox_2_and_516
      ^ Encrypt_Top_sbox_2_and_652;
  assign xor_cse_189 = state_2_11_1_lpi_4 ^ state_0_11_lpi_6 ^ state_3_11_lpi_3 ^
      state_1_1_31_0_lpi_4_11;
  assign xor_cse_190 = Encrypt_Top_sbox_1_and_1_cse_11_sva_1 ^ Encrypt_Top_sbox_1_and_cse_11_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1 ^ state_0_47_lpi_6;
  assign xor_cse_188 = xor_cse_189 ^ xor_cse_84 ^ xor_cse_190 ^ Encrypt_Top_sbox_1_and_1_cse_47_sva_1;
  assign xor_cse_192 = state_1_1_63_32_lpi_4_15 ^ (state_4_4_47_lpi_3 & state_1_1_63_32_lpi_4_15)
      ^ state_3_47_lpi_3 ^ (state_1_1_63_32_lpi_4_15 & state_0_47_lpi_6);
  assign ciphertext_47_sva_mx0w2 = xor_cse_188 ^ xor_cse_192 ^ xor_cse_88 ^ plaintext_63_32_sva_15
      ^ state_2_47_1_lpi_4;
  assign xor_cse_194 = xor_cse_119 ^ Encrypt_Top_sbox_2_and_566 ^ Encrypt_Top_sbox_2_and_564
      ^ Encrypt_Top_sbox_2_and_644;
  assign xor_cse_196 = state_1_1_31_0_lpi_4_0 ^ state_3_0_lpi_3 ^ state_0_0_lpi_6
      ^ state_4_4_0_lpi_3;
  assign xor_cse_197 = state_2_0_1_lpi_4 ^ Encrypt_Top_sbox_2_and_520 ^ Encrypt_Top_sbox_2_and_522
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0]);
  assign xor_cse_195 = xor_cse_196 ^ xor_cse_197 ^ Encrypt_Top_sbox_2_and_646 ^ state_1_1_63_32_lpi_4_20;
  assign xor_cse_201 = state_1_1_63_32_lpi_4_16 ^ (state_4_4_48_lpi_3 & state_1_1_63_32_lpi_4_16)
      ^ state_3_48_lpi_3 ^ (state_1_1_63_32_lpi_4_16 & state_0_48_lpi_6);
  assign xor_cse_202 = Encrypt_Top_sbox_1_and_1_cse_12_sva_1 ^ Encrypt_Top_sbox_1_and_cse_12_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_12_sva_1 ^ state_0_48_lpi_6;
  assign xor_cse_200 = Encrypt_Top_sbox_1_and_1_cse_48_sva_1 ^ state_2_48_1_lpi_4
      ^ xor_cse_201 ^ xor_cse_202;
  assign xor_cse_204 = state_2_12_1_lpi_4 ^ state_0_12_lpi_6 ^ state_3_12_lpi_3 ^
      state_1_1_31_0_lpi_4_12;
  assign ciphertext_48_sva_mx0w2 = xor_cse_200 ^ plaintext_63_32_sva_16 ^ xor_cse_204
      ^ xor_cse_102 ^ xor_cse_103;
  assign xor_cse_206 = state_1_1_31_0_lpi_4_1 ^ state_3_1_lpi_3 ^ state_0_1_lpi_6
      ^ state_4_4_1_lpi_3;
  assign xor_cse_207 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1])
      ^ Encrypt_Top_sbox_2_and_528 ^ Encrypt_Top_sbox_2_and_530;
  assign xor_cse_205 = xor_cse_206 ^ xor_cse_207 ^ Encrypt_Top_sbox_2_and_558 ^ state_1_1_63_32_lpi_4_30;
  assign xor_cse_209 = state_1_1_63_32_lpi_4_21 ^ Encrypt_Top_sbox_2_and_636 ^ Encrypt_Top_sbox_2_and_638
      ^ Encrypt_Top_sbox_2_and_556;
  assign xor_cse_211 = state_2_13_1_lpi_4 ^ state_0_13_lpi_6 ^ state_3_13_lpi_3 ^
      state_1_1_31_0_lpi_4_13;
  assign xor_cse_210 = xor_cse_211 ^ state_0_49_lpi_6 ^ xor_cse_111 ^ Encrypt_Top_sbox_1_and_1_cse_13_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_13_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1
      ^ state_2_49_1_lpi_4;
  assign xor_cse_214 = state_1_1_63_32_lpi_4_17 ^ (state_4_4_49_lpi_3 & state_1_1_63_32_lpi_4_17)
      ^ state_3_49_lpi_3 ^ (state_1_1_63_32_lpi_4_17 & state_0_49_lpi_6);
  assign ciphertext_49_sva_mx0w2 = xor_cse_210 ^ xor_cse_214 ^ xor_cse_116 ^ plaintext_63_32_sva_17
      ^ Encrypt_Top_sbox_1_and_1_cse_49_sva_1;
  assign xor_cse_217 = state_1_1_31_0_lpi_4_2 ^ state_3_2_lpi_3 ^ state_0_2_lpi_6
      ^ state_4_4_2_lpi_3;
  assign xor_cse_218 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ Encrypt_Top_sbox_2_and_536 ^ Encrypt_Top_sbox_2_and_538;
  assign xor_cse_221 = state_2_14_1_lpi_4 ^ state_0_14_lpi_6 ^ state_3_14_lpi_3 ^
      state_1_1_31_0_lpi_4_14;
  assign xor_cse_222 = Encrypt_Top_sbox_1_and_1_cse_14_sva_1 ^ Encrypt_Top_sbox_1_and_cse_14_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1 ^ state_0_50_lpi_6;
  assign xor_cse_220 = xor_cse_221 ^ xor_cse_124 ^ xor_cse_222 ^ Encrypt_Top_sbox_1_and_1_cse_50_sva_1;
  assign xor_cse_224 = state_1_1_63_32_lpi_4_18 ^ (state_4_4_50_lpi_3 & state_1_1_63_32_lpi_4_18)
      ^ state_3_50_lpi_3 ^ (state_1_1_63_32_lpi_4_18 & state_0_50_lpi_6);
  assign ciphertext_50_sva_mx0w2 = xor_cse_220 ^ xor_cse_224 ^ xor_cse_125 ^ plaintext_63_32_sva_18
      ^ state_2_50_1_lpi_4;
  assign xor_cse_226 = xor_cse_24 ^ Encrypt_Top_sbox_2_and_622 ^ Encrypt_Top_sbox_2_and_620
      ^ state_1_1_63_32_lpi_4_23;
  assign xor_cse_228 = state_1_1_31_0_lpi_4_3 ^ state_3_3_lpi_3 ^ state_0_3_lpi_6
      ^ state_4_4_3_lpi_3;
  assign xor_cse_229 = state_2_3_1_lpi_4 ^ Encrypt_Top_sbox_2_and_544 ^ Encrypt_Top_sbox_2_and_546
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3]);
  assign xor_cse_231 = state_2_15_1_lpi_4 ^ state_0_15_lpi_6 ^ state_3_15_lpi_3 ^
      state_1_1_31_0_lpi_4_15;
  assign xor_cse_230 = xor_cse_136 ^ state_0_51_lpi_6 ^ xor_cse_231 ^ Encrypt_Top_sbox_1_and_1_cse_15_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_15_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1
      ^ state_2_51_1_lpi_4;
  assign ciphertext_51_sva_mx0w2 = xor_cse_230 ^ xor_cse_1 ^ xor_cse_137 ^ plaintext_63_32_sva_19
      ^ Encrypt_Top_sbox_1_and_1_cse_51_sva_1;
  assign xor_cse_236 = Encrypt_Top_sbox_2_and_534 ^ Encrypt_Top_sbox_2_and_532 ^
      Encrypt_Top_sbox_2_and_612 ^ Encrypt_Top_sbox_2_and_614;
  assign xor_cse_235 = xor_cse_37 ^ xor_cse_164 ^ xor_cse_236 ^ state_1_1_63_32_lpi_4_24;
  assign xor_cse_238 = state_1_1_31_0_lpi_4_4 ^ state_3_4_lpi_3 ^ state_0_4_lpi_6
      ^ state_4_4_4_lpi_3;
  assign xor_cse_239 = state_2_4_1_lpi_4 ^ Encrypt_Top_sbox_2_and_552 ^ Encrypt_Top_sbox_2_and_554
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4]);
  assign xor_cse_242 = state_2_16_1_lpi_4 ^ state_0_16_lpi_6 ^ state_3_16_lpi_3 ^
      state_1_1_31_0_lpi_4_16;
  assign xor_cse_241 = xor_cse_242 ^ state_0_52_lpi_6 ^ xor_cse_148 ^ Encrypt_Top_sbox_1_and_1_cse_16_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_16_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1
      ^ state_2_52_1_lpi_4;
  assign ciphertext_52_sva_mx0w2 = xor_cse_241 ^ xor_cse_15 ^ xor_cse_149 ^ plaintext_63_32_sva_20
      ^ Encrypt_Top_sbox_1_and_1_cse_52_sva_1;
  assign xor_cse_246 = xor_cse_174 ^ Encrypt_Top_sbox_2_and_526 ^ Encrypt_Top_sbox_2_and_524
      ^ Encrypt_Top_sbox_2_and_604;
  assign xor_cse_248 = state_1_1_31_0_lpi_4_5 ^ state_3_5_lpi_3 ^ state_0_5_lpi_6
      ^ state_4_4_5_lpi_3;
  assign xor_cse_249 = state_2_5_1_lpi_4 ^ Encrypt_Top_sbox_2_and_560 ^ Encrypt_Top_sbox_2_and_562
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5]);
  assign xor_cse_252 = state_2_17_1_lpi_4 ^ state_0_17_lpi_6 ^ state_3_17_lpi_3 ^
      state_1_1_31_0_lpi_4_17;
  assign xor_cse_251 = xor_cse_252 ^ Encrypt_Top_sbox_1_and_1_cse_17_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_17_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_17_sva_1;
  assign xor_cse_254 = state_2_53_1_lpi_4 ^ state_0_53_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_53_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_8_sva_1;
  assign ciphertext_53_sva_mx0w2 = xor_cse_251 ^ xor_cse_29 ^ xor_cse_159 ^ xor_cse_254
      ^ plaintext_63_32_sva_21 ^ state_2_8_1_lpi_4 ^ state_0_8_lpi_6;
  assign xor_cse_256 = xor_cse_65 ^ Encrypt_Top_sbox_2_and_598 ^ Encrypt_Top_sbox_2_and_516
      ^ Encrypt_Top_sbox_2_and_518;
  assign xor_cse_258 = state_1_1_31_0_lpi_4_6 ^ state_3_6_lpi_3 ^ state_0_6_lpi_6
      ^ state_4_4_6_lpi_3;
  assign xor_cse_257 = xor_cse_185 ^ xor_cse_258 ^ Encrypt_Top_sbox_2_and_596 ^ state_1_1_63_32_lpi_4_26;
  assign xor_cse_260 = state_2_6_1_lpi_4 ^ Encrypt_Top_sbox_2_and_568 ^ Encrypt_Top_sbox_2_and_570
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6]);
  assign xor_cse_263 = state_2_18_1_lpi_4 ^ state_0_18_lpi_6 ^ state_3_18_lpi_3 ^
      state_1_1_31_0_lpi_4_18;
  assign xor_cse_262 = state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ state_0_54_lpi_6 ^ xor_cse_263;
  assign xor_cse_265 = Encrypt_Top_sbox_1_and_1_cse_18_sva_1 ^ Encrypt_Top_sbox_1_and_cse_18_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1 ^ state_2_54_1_lpi_4;
  assign ciphertext_54_sva_mx0w2 = xor_cse_262 ^ xor_cse_44 ^ xor_cse_170 ^ xor_cse_265
      ^ plaintext_63_32_sva_22 ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_9_sva_1;
  assign xor_cse_268 = state_1_1_31_0_lpi_4_7 ^ state_3_7_lpi_3 ^ state_0_7_lpi_6
      ^ state_4_4_7_lpi_3;
  assign xor_cse_267 = xor_cse_79 ^ Encrypt_Top_sbox_2_and_588 ^ Encrypt_Top_sbox_2_and_590
      ^ xor_cse_268;
  assign xor_cse_270 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7])
      ^ Encrypt_Top_sbox_2_and_576 ^ Encrypt_Top_sbox_2_and_578;
  assign xor_cse_272 = xor_cse_178 ^ Encrypt_Top_sbox_1_and_cse_10_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_10_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_10_sva_1;
  assign xor_cse_274 = state_2_19_1_lpi_4 ^ state_0_19_lpi_6 ^ state_3_19_lpi_3 ^
      state_1_1_31_0_lpi_4_19;
  assign xor_cse_275 = Encrypt_Top_sbox_1_and_1_cse_19_sva_1 ^ Encrypt_Top_sbox_1_and_cse_19_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1 ^ state_2_55_1_lpi_4;
  assign ciphertext_55_sva_mx0w2 = xor_cse_272 ^ xor_cse_274 ^ xor_cse_57 ^ xor_cse_275
      ^ plaintext_63_32_sva_23 ^ Encrypt_Top_sbox_1_and_1_cse_55_sva_1 ^ state_0_55_lpi_6;
  assign xor_cse_278 = state_2_8_1_lpi_4 ^ state_0_8_lpi_6 ^ state_3_8_lpi_3 ^ state_4_4_8_lpi_3;
  assign xor_cse_277 = xor_cse_278 ^ Encrypt_Top_sbox_2_and_586 ^ Encrypt_Top_sbox_2_and_584
      ^ state_1_1_63_32_lpi_4_8;
  assign xor_cse_280 = xor_cse_189 ^ Encrypt_Top_sbox_1_and_cse_11_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_11_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1;
  assign xor_cse_282 = state_2_20_1_lpi_4 ^ state_0_20_lpi_6 ^ state_3_20_lpi_3 ^
      state_1_1_31_0_lpi_4_20;
  assign xor_cse_283 = Encrypt_Top_sbox_1_and_1_cse_20_sva_1 ^ Encrypt_Top_sbox_1_and_cse_20_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1 ^ state_2_56_1_lpi_4;
  assign ciphertext_56_sva_mx0w2 = xor_cse_280 ^ xor_cse_282 ^ xor_cse_73 ^ xor_cse_283
      ^ plaintext_63_32_sva_24 ^ Encrypt_Top_sbox_1_and_1_cse_56_sva_1 ^ state_0_56_lpi_6;
  assign xor_cse_286 = state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ state_3_9_lpi_3 ^ state_4_4_9_lpi_3;
  assign xor_cse_285 = xor_cse_286 ^ Encrypt_Top_sbox_2_and_592 ^ Encrypt_Top_sbox_2_and_594
      ^ state_1_1_63_32_lpi_4_9;
  assign xor_cse_288 = xor_cse_204 ^ Encrypt_Top_sbox_1_and_cse_12_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_12_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_12_sva_1;
  assign xor_cse_290 = state_2_21_1_lpi_4 ^ state_0_21_lpi_6 ^ state_3_21_lpi_3 ^
      state_1_1_31_0_lpi_4_21;
  assign xor_cse_291 = Encrypt_Top_sbox_1_and_1_cse_21_sva_1 ^ Encrypt_Top_sbox_1_and_cse_21_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1 ^ state_2_57_1_lpi_4;
  assign ciphertext_57_sva_mx0w2 = xor_cse_288 ^ xor_cse_290 ^ xor_cse_85 ^ xor_cse_291
      ^ plaintext_63_32_sva_25 ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1 ^ state_0_57_lpi_6;
  assign xor_cse_293 = xor_cse_119 ^ Encrypt_Top_sbox_2_and_566 ^ xor_cse_178 ^ state_4_4_10_lpi_3
      ^ Encrypt_Top_sbox_2_and_600 ^ Encrypt_Top_sbox_2_and_602 ^ Encrypt_Top_sbox_2_and_564;
  assign xor_cse_297 = xor_cse_211 ^ Encrypt_Top_sbox_1_and_cse_13_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_13_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1;
  assign xor_cse_299 = state_2_22_1_lpi_4 ^ state_0_22_lpi_6 ^ state_3_22_lpi_3 ^
      state_1_1_31_0_lpi_4_22;
  assign xor_cse_300 = Encrypt_Top_sbox_1_and_cse_22_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_22_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_22_sva_1 ^ state_2_58_1_lpi_4;
  assign ciphertext_58_sva_mx0w2 = xor_cse_297 ^ xor_cse_299 ^ xor_cse_100 ^ xor_cse_300
      ^ plaintext_63_32_sva_26 ^ Encrypt_Top_sbox_1_and_1_cse_58_sva_1 ^ state_0_58_lpi_6;
  assign xor_cse_302 = xor_cse_189 ^ Encrypt_Top_sbox_2_and_558 ^ xor_cse_132 ^ state_4_4_11_lpi_3
      ^ Encrypt_Top_sbox_2_and_608 ^ Encrypt_Top_sbox_2_and_610 ^ Encrypt_Top_sbox_2_and_556;
  assign xor_cse_306 = xor_cse_221 ^ Encrypt_Top_sbox_1_and_cse_14_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_14_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1;
  assign xor_cse_308 = state_2_23_1_lpi_4 ^ state_0_23_lpi_6 ^ state_3_23_lpi_3 ^
      state_1_1_31_0_lpi_4_23;
  assign xor_cse_309 = Encrypt_Top_sbox_1_and_1_cse_23_sva_1 ^ Encrypt_Top_sbox_1_and_cse_23_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1 ^ state_0_59_lpi_6;
  assign ciphertext_59_sva_mx0w2 = xor_cse_306 ^ xor_cse_308 ^ xor_cse_115 ^ xor_cse_309
      ^ plaintext_63_32_sva_27 ^ Encrypt_Top_sbox_1_and_1_cse_59_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1;
  assign xor_cse_311 = xor_cse_204 ^ Encrypt_Top_sbox_2_and_550 ^ xor_cse_142 ^ state_4_4_12_lpi_3
      ^ Encrypt_Top_sbox_2_and_616 ^ Encrypt_Top_sbox_2_and_618 ^ Encrypt_Top_sbox_2_and_548;
  assign xor_cse_316 = state_2_24_1_lpi_4 ^ state_0_24_lpi_6 ^ state_3_24_lpi_3 ^
      state_1_1_31_0_lpi_4_24;
  assign xor_cse_315 = xor_cse_231 ^ Encrypt_Top_sbox_1_and_1_cse_15_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1
      ^ xor_cse_316;
  assign xor_cse_318 = Encrypt_Top_sbox_1_and_cse_24_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_24_sva_1 ^ Encrypt_Top_sbox_1_and_cse_15_sva_1;
  assign ciphertext_60_sva_mx0w2 = xor_cse_315 ^ xor_cse_3 ^ xor_cse_318 ^ plaintext_63_32_sva_28
      ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_60_sva_1
      ^ state_1_1_63_32_lpi_4_28;
  assign xor_cse_320 = xor_cse_154 ^ Encrypt_Top_sbox_2_and_542 ^ xor_cse_211 ^ state_4_4_13_lpi_3
      ^ Encrypt_Top_sbox_2_and_624 ^ Encrypt_Top_sbox_2_and_626 ^ Encrypt_Top_sbox_2_and_540;
  assign xor_cse_325 = state_2_25_1_lpi_4 ^ state_0_25_lpi_6 ^ state_3_25_lpi_3 ^
      state_1_1_31_0_lpi_4_25;
  assign xor_cse_324 = Encrypt_Top_sbox_2_and_2_cse_25_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_25_sva_1
      ^ xor_cse_325 ^ xor_cse_242;
  assign xor_cse_327 = Encrypt_Top_sbox_1_and_1_cse_16_sva_1 ^ Encrypt_Top_sbox_1_and_cse_16_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1 ^ Encrypt_Top_sbox_1_and_cse_25_sva_1;
  assign ciphertext_61_sva_mx0w2 = xor_cse_324 ^ xor_cse_17 ^ xor_cse_327 ^ plaintext_63_32_sva_29
      ^ Encrypt_Top_sbox_1_and_1_cse_61_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_61_sva_1
      ^ state_1_1_63_32_lpi_4_29;
  assign xor_cse_329 = xor_cse_268 ^ Encrypt_Top_sbox_2_and_534 ^ xor_cse_164 ^ xor_cse_221;
  assign xor_cse_331 = state_4_4_14_lpi_3 ^ Encrypt_Top_sbox_2_and_632 ^ Encrypt_Top_sbox_2_and_634
      ^ Encrypt_Top_sbox_2_and_532;
  assign xor_cse_334 = state_2_26_1_lpi_4 ^ state_0_26_lpi_6 ^ state_3_26_lpi_3 ^
      state_1_1_31_0_lpi_4_26;
  assign xor_cse_333 = xor_cse_252 ^ Encrypt_Top_sbox_1_and_1_cse_17_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_17_sva_1
      ^ xor_cse_334;
  assign xor_cse_336 = Encrypt_Top_sbox_1_and_cse_26_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_26_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_26_sva_1 ^ Encrypt_Top_sbox_1_and_cse_17_sva_1;
  assign ciphertext_62_sva_mx0w2 = xor_cse_333 ^ xor_cse_28 ^ xor_cse_336 ^ plaintext_63_32_sva_30
      ^ Encrypt_Top_sbox_1_and_1_cse_62_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_62_sva_1
      ^ state_1_1_63_32_lpi_4_30;
  assign xor_cse_339 = state_4_4_15_lpi_3 ^ Encrypt_Top_sbox_2_and_640 ^ Encrypt_Top_sbox_2_and_642
      ^ Encrypt_Top_sbox_2_and_524;
  assign xor_cse_341 = xor_cse_263 ^ Encrypt_Top_sbox_1_and_cse_18_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_18_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1;
  assign xor_cse_343 = state_2_27_1_lpi_4 ^ state_0_27_lpi_6 ^ state_3_27_lpi_3 ^
      state_1_1_31_0_lpi_4_27;
  assign xor_cse_344 = Encrypt_Top_sbox_1_and_cse_27_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_27_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_27_sva_1 ^ state_2_63_1_lpi_4;
  assign ciphertext_63_sva_mx0w2 = xor_cse_341 ^ xor_cse_343 ^ xor_cse_42 ^ xor_cse_344
      ^ plaintext_63_32_sva_31 ^ Encrypt_Top_sbox_1_and_1_cse_63_sva_1 ^ state_0_63_lpi_6;
  assign xor_cse_347 = state_4_4_16_lpi_3 ^ Encrypt_Top_sbox_2_and_648 ^ Encrypt_Top_sbox_2_and_650
      ^ Encrypt_Top_sbox_2_and_516;
  assign xor_cse_350 = plaintext_31_0_sva_19 ^ (state_4_3_31_0_sva_19 & plaintext_31_0_sva_19)
      ^ state_3_3_31_0_sva_19 ^ (plaintext_31_0_sva_19 & state_0_19_lpi_6);
  assign xor_cse_349 = state_2_19_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_19_sva_1 ^
      state_0_19_lpi_6 ^ xor_cse_350;
  assign xor_cse_352 = state_2_0_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0])
      ^ state_0_0_lpi_6 ^ state_3_3_31_0_sva_0;
  assign xor_cse_351 = xor_cse_352 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_0 ^ Encrypt_Top_sbox_and_1_cse_0_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_0_sva_1;
  assign xor_cse_354 = plaintext_31_0_sva_28 ^ (state_4_3_31_0_sva_28 & plaintext_31_0_sva_28)
      ^ state_3_3_31_0_sva_28 ^ (plaintext_31_0_sva_28 & state_0_28_lpi_6);
  assign xor_cse_357 = state_2_28_1_lpi_4 ^ state_0_28_lpi_6 ^ state_3_28_lpi_3 ^
      state_1_1_31_0_lpi_4_28;
  assign xor_cse_356 = xor_cse_357 ^ Encrypt_Top_sbox_1_and_cse_28_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_28_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_28_sva_1;
  assign xor_cse_358 = xor_cse_274 ^ Encrypt_Top_sbox_1_and_cse_19_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_19_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1;
  assign xor_cse_359 = state_2_0_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_0_sva_1 ^
      (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]) ^ state_0_0_lpi_6;
  assign xor_cse_360 = state_2_0_1_lpi_4 ^ state_0_0_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_0_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0]);
  assign xor_cse_362 = plaintext_31_0_sva_20 ^ (state_4_3_31_0_sva_20 & plaintext_31_0_sva_20)
      ^ state_3_3_31_0_sva_20 ^ (plaintext_31_0_sva_20 & state_0_20_lpi_6);
  assign xor_cse_361 = state_2_20_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_20_sva_1 ^
      state_0_20_lpi_6 ^ xor_cse_362;
  assign xor_cse_364 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1])
      ^ state_0_1_lpi_6 ^ state_3_3_31_0_sva_1;
  assign xor_cse_363 = xor_cse_364 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_1 ^ Encrypt_Top_sbox_and_1_cse_1_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_1_sva_1;
  assign xor_cse_366 = plaintext_31_0_sva_29 ^ (state_4_3_31_0_sva_29 & plaintext_31_0_sva_29)
      ^ state_3_3_31_0_sva_29 ^ (plaintext_31_0_sva_29 & state_0_29_lpi_6);
  assign xor_cse_369 = state_2_29_1_lpi_4 ^ state_0_29_lpi_6 ^ state_3_29_lpi_3 ^
      state_1_1_31_0_lpi_4_29;
  assign xor_cse_368 = xor_cse_369 ^ Encrypt_Top_sbox_1_and_cse_29_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_29_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_29_sva_1;
  assign xor_cse_370 = xor_cse_282 ^ Encrypt_Top_sbox_1_and_cse_20_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_20_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1;
  assign xor_cse_373 = state_2_1_1_lpi_4 ^ state_0_1_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_1_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1]);
  assign xor_cse_375 = plaintext_31_0_sva_21 ^ (state_4_3_31_0_sva_21 & plaintext_31_0_sva_21)
      ^ state_3_3_31_0_sva_21 ^ (plaintext_31_0_sva_21 & state_0_21_lpi_6);
  assign xor_cse_374 = state_2_21_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_21_sva_1 ^
      state_0_21_lpi_6 ^ xor_cse_375;
  assign xor_cse_377 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ state_0_2_lpi_6 ^ state_3_3_31_0_sva_2;
  assign xor_cse_376 = xor_cse_377 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_2 ^ Encrypt_Top_sbox_and_1_cse_2_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_2_sva_1;
  assign xor_cse_379 = plaintext_31_0_sva_30 ^ (state_4_3_31_0_sva_30 & plaintext_31_0_sva_30)
      ^ state_3_3_31_0_sva_30 ^ (plaintext_31_0_sva_30 & state_0_30_lpi_6);
  assign xor_cse_381 = Encrypt_Top_sbox_1_and_cse_30_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_30_sva_1 ^ Encrypt_Top_sbox_1_and_cse_21_sva_1;
  assign xor_cse_382 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2])
      ^ Encrypt_Top_sbox_1_and_1_cse_2_sva_1 ^ state_0_2_lpi_6;
  assign xor_cse_384 = state_2_30_1_lpi_4 ^ state_0_30_lpi_6 ^ state_3_30_lpi_3 ^
      state_1_1_31_0_lpi_4_30;
  assign xor_cse_383 = xor_cse_290 ^ Encrypt_Top_sbox_1_and_1_cse_21_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1
      ^ xor_cse_384;
  assign xor_cse_385 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ Encrypt_Top_sbox_3_and_1_cse_2_sva_1 ^ state_0_2_lpi_6;
  assign xor_cse_387 = plaintext_31_0_sva_22 ^ (state_4_3_31_0_sva_22 & plaintext_31_0_sva_22)
      ^ state_3_3_31_0_sva_22 ^ (plaintext_31_0_sva_22 & state_0_22_lpi_6);
  assign xor_cse_386 = state_2_22_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_22_sva_1 ^
      state_0_22_lpi_6 ^ xor_cse_387;
  assign xor_cse_389 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ state_0_3_lpi_6 ^ state_3_3_31_0_sva_3;
  assign xor_cse_390 = plaintext_31_0_sva_31 ^ (state_4_3_31_0_sva_31 & plaintext_31_0_sva_31)
      ^ state_3_3_31_0_sva_31 ^ (plaintext_31_0_sva_31 & state_0_31_lpi_6);
  assign xor_cse_394 = state_2_31_1_lpi_4 ^ state_0_31_lpi_6 ^ state_3_31_lpi_3 ^
      state_1_1_31_0_lpi_4_31;
  assign xor_cse_393 = xor_cse_394 ^ Encrypt_Top_sbox_1_and_cse_31_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_31_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_31_sva_1;
  assign xor_cse_395 = xor_cse_299 ^ Encrypt_Top_sbox_1_and_cse_22_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_22_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_22_sva_1;
  assign xor_cse_401 = state_2_32_1_lpi_4 ^ state_0_32_lpi_6 ^ plaintext_63_32_sva_0
      ^ state_3_3_63_32_sva_0;
  assign xor_cse_400 = xor_cse_401 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_0 ^ Encrypt_Top_sbox_and_1_cse_32_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_32_sva_1;
  assign xor_cse_403 = plaintext_31_0_sva_23 ^ (state_4_3_31_0_sva_23 & plaintext_31_0_sva_23)
      ^ state_3_3_31_0_sva_23 ^ (plaintext_31_0_sva_23 & state_0_23_lpi_6);
  assign xor_cse_402 = state_2_23_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_23_sva_1 ^
      state_0_23_lpi_6 ^ xor_cse_403;
  assign xor_cse_405 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4])
      ^ state_0_4_lpi_6 ^ state_3_3_31_0_sva_4;
  assign xor_cse_407 = xor_cse_308 ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1 ^ xor_cse_111
      ^ state_2_32_1_lpi_4 ^ state_0_32_lpi_6 ^ Encrypt_Top_sbox_1_and_cse_23_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_23_sva_1;
  assign state_0_4_sva_4_mx0w4 = Encrypt_Top_sbox_1_and_1_cse_32_sva_1 ^ xor_cse_4
      ^ xor_cse_116 ^ xor_cse_407;
  assign xor_cse_412 = state_1_1_31_0_lpi_4_8 ^ (state_4_4_32_lpi_3 & state_1_1_31_0_lpi_4_8)
      ^ state_3_32_lpi_3 ^ (state_1_1_31_0_lpi_4_8 & state_0_32_lpi_6);
  assign xor_cse_415 = plaintext_31_0_sva_24 ^ (state_4_3_31_0_sva_24 & plaintext_31_0_sva_24)
      ^ state_3_3_31_0_sva_24 ^ (plaintext_31_0_sva_24 & state_0_24_lpi_6);
  assign xor_cse_414 = state_2_24_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_24_sva_1 ^
      state_0_24_lpi_6 ^ xor_cse_415;
  assign xor_cse_417 = state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5])
      ^ state_0_5_lpi_6 ^ state_3_3_31_0_sva_5;
  assign xor_cse_416 = xor_cse_417 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_5 ^ Encrypt_Top_sbox_and_1_cse_5_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_5_sva_1;
  assign xor_cse_419 = state_2_33_1_lpi_4 ^ state_0_33_lpi_6 ^ plaintext_63_32_sva_1
      ^ state_3_3_63_32_sva_1;
  assign xor_cse_421 = xor_cse_124 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1 ^ xor_cse_316
      ^ state_2_33_1_lpi_4 ^ state_0_33_lpi_6 ^ Encrypt_Top_sbox_1_and_cse_24_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_24_sva_1;
  assign state_0_5_sva_4_mx0w4 = Encrypt_Top_sbox_1_and_1_cse_33_sva_1 ^ xor_cse_125
      ^ xor_cse_18 ^ xor_cse_421;
  assign xor_cse_425 = state_1_1_31_0_lpi_4_9 ^ (state_4_4_33_lpi_3 & state_1_1_31_0_lpi_4_9)
      ^ state_3_33_lpi_3 ^ (state_1_1_31_0_lpi_4_9 & state_0_33_lpi_6);
  assign xor_cse_426 = state_2_5_1_lpi_4 ^ state_0_5_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_5_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5]);
  assign xor_cse_428 = plaintext_31_0_sva_25 ^ (state_4_3_31_0_sva_25 & plaintext_31_0_sva_25)
      ^ state_3_3_31_0_sva_25 ^ (plaintext_31_0_sva_25 & state_0_25_lpi_6);
  assign xor_cse_427 = state_2_25_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_25_sva_1 ^
      state_0_25_lpi_6 ^ xor_cse_428;
  assign xor_cse_430 = state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6])
      ^ state_0_6_lpi_6 ^ state_3_3_31_0_sva_6;
  assign xor_cse_431 = state_2_34_1_lpi_4 ^ state_0_34_lpi_6 ^ plaintext_63_32_sva_2
      ^ state_3_3_63_32_sva_2;
  assign xor_cse_434 = state_2_34_1_lpi_4 ^ state_0_34_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_25_sva_1;
  assign xor_cse_435 = state_2_6_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_6_sva_1 ^
      (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]) ^ state_0_6_lpi_6;
  assign xor_cse_436 = Encrypt_Top_sbox_1_and_1_cse_25_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1;
  assign state_0_6_sva_4_mx0w4 = xor_cse_325 ^ xor_cse_136 ^ xor_cse_30 ^ xor_cse_137
      ^ xor_cse_434 ^ xor_cse_436;
  assign xor_cse_439 = state_1_1_63_32_lpi_4_0 ^ (state_4_4_34_lpi_3 & state_1_1_63_32_lpi_4_0)
      ^ state_3_34_lpi_3 ^ (state_1_1_63_32_lpi_4_0 & state_0_34_lpi_6);
  assign xor_cse_438 = state_2_34_1_lpi_4 ^ state_0_34_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_34_sva_1
      ^ xor_cse_439;
  assign xor_cse_441 = state_2_6_1_lpi_4 ^ state_0_6_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_6_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6]);
  assign xor_cse_444 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7])
      ^ state_0_7_lpi_6 ^ state_3_3_31_0_sva_7;
  assign xor_cse_443 = xor_cse_444 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_7 ^ Encrypt_Top_sbox_and_1_cse_7_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_7_sva_1;
  assign xor_cse_446 = state_2_35_1_lpi_4 ^ state_0_35_lpi_6 ^ plaintext_63_32_sva_3
      ^ state_3_3_63_32_sva_3;
  assign xor_cse_445 = xor_cse_446 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_3 ^ Encrypt_Top_sbox_and_1_cse_35_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_35_sva_1;
  assign xor_cse_448 = plaintext_31_0_sva_26 ^ (state_4_3_31_0_sva_26 & plaintext_31_0_sva_26)
      ^ state_3_3_31_0_sva_26 ^ (plaintext_31_0_sva_26 & state_0_26_lpi_6);
  assign xor_cse_450 = xor_cse_334 ^ Encrypt_Top_sbox_1_and_cse_26_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_26_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_26_sva_1;
  assign xor_cse_452 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7])
      ^ Encrypt_Top_sbox_1_and_1_cse_7_sva_1 ^ state_0_7_lpi_6;
  assign xor_cse_453 = Encrypt_Top_sbox_1_and_1_cse_35_sva_1 ^ state_2_35_1_lpi_4
      ^ state_0_35_lpi_6;
  assign state_0_7_sva_4_mx0w4 = xor_cse_450 ^ xor_cse_148 ^ xor_cse_46 ^ xor_cse_149
      ^ xor_cse_453;
  assign xor_cse_456 = state_2_7_1_lpi_4 ^ state_0_7_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_7_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7]);
  assign xor_cse_458 = state_1_1_63_32_lpi_4_1 ^ (state_4_4_35_lpi_3 & state_1_1_63_32_lpi_4_1)
      ^ state_3_35_lpi_3 ^ (state_1_1_63_32_lpi_4_1 & state_0_35_lpi_6);
  assign xor_cse_457 = state_2_35_1_lpi_4 ^ state_0_35_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_35_sva_1
      ^ xor_cse_458;
  assign xor_cse_459 = state_2_16_1_lpi_4 ^ (state_4_3_31_0_sva_16 & state_3_3_31_0_sva_16)
      ^ state_4_3_31_0_sva_16 ^ plaintext_31_0_sva_16;
  assign xor_cse_462 = state_4_3_31_0_sva_10 & state_3_3_31_0_sva_10;
  assign xor_cse_461 = xor_cse_462 ^ state_4_3_31_0_sva_10 ^ state_2_10_1_lpi_4 ^
      plaintext_31_0_sva_10;
  assign xor_cse_464 = state_4_3_31_0_sva_11 & state_3_3_31_0_sva_11;
  assign xor_cse_463 = xor_cse_464 ^ state_4_3_31_0_sva_11 ^ state_2_11_1_lpi_4 ^
      plaintext_31_0_sva_11;
  assign xor_cse_465 = state_4_4_10_lpi_3 ^ state_1_1_31_0_lpi_4_10 ^ (state_4_4_10_lpi_3
      & state_3_10_lpi_3) ^ state_2_10_1_lpi_4;
  assign xor_cse_466 = state_2_11_1_lpi_4 ^ (state_4_4_11_lpi_3 & state_3_11_lpi_3)
      ^ state_4_4_11_lpi_3 ^ state_1_1_31_0_lpi_4_11;
  assign xor_cse_467 = Encrypt_Top_sbox_1_and_784 ^ state_4_4_16_lpi_3 ^ state_2_16_1_lpi_4
      ^ state_1_1_31_0_lpi_4_16;
  assign xor_cse_468 = state_4_4_23_lpi_3 ^ state_1_1_31_0_lpi_4_23 ^ Encrypt_Top_sbox_1_and_cse_23_sva_1
      ^ state_3_23_lpi_3;
  assign xor_cse_469 = state_4_4_16_lpi_3 ^ state_1_1_31_0_lpi_4_16 ^ Encrypt_Top_sbox_1_and_cse_16_sva_1
      ^ state_3_16_lpi_3;
  assign xor_cse_470 = state_1_1_63_32_lpi_4_3 ^ (state_4_4_57_lpi_3 & state_1_1_63_32_lpi_4_3)
      ^ state_3_57_lpi_3 ^ (state_1_1_63_32_lpi_4_3 & state_0_57_lpi_6);
  assign xor_cse_471 = Encrypt_Top_sbox_2_and_2_cse_16_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1
      ^ state_4_4_57_lpi_3;
  assign state_4_16_sva_2_mx0w4 = xor_cse_468 ^ xor_cse_469 ^ xor_cse_470 ^ xor_cse_471;
  assign xor_cse_472 = state_4_3_31_0_sva_17 ^ (state_4_3_31_0_sva_17 & state_3_3_31_0_sva_17)
      ^ state_2_17_1_lpi_4 ^ plaintext_31_0_sva_17;
  assign xor_cse_476 = state_4_3_31_0_sva_12 & state_3_3_31_0_sva_12;
  assign xor_cse_475 = xor_cse_476 ^ state_4_3_31_0_sva_12 ^ state_2_12_1_lpi_4 ^
      plaintext_31_0_sva_12;
  assign xor_cse_477 = state_2_12_1_lpi_4 ^ (state_4_4_12_lpi_3 & state_3_12_lpi_3)
      ^ state_4_4_12_lpi_3 ^ state_1_1_31_0_lpi_4_12;
  assign xor_cse_479 = state_4_4_17_lpi_3 ^ state_1_1_31_0_lpi_4_17 ^ Encrypt_Top_sbox_1_and_cse_17_sva_1
      ^ state_3_17_lpi_3;
  assign xor_cse_480 = state_1_1_63_32_lpi_4_30 ^ (state_4_4_58_lpi_3 & state_1_1_63_32_lpi_4_30)
      ^ state_3_58_lpi_3 ^ (state_1_1_63_32_lpi_4_30 & state_0_58_lpi_6);
  assign xor_cse_481 = state_4_4_24_lpi_3 ^ state_1_1_31_0_lpi_4_24 ^ Encrypt_Top_sbox_1_and_cse_24_sva_1
      ^ state_3_24_lpi_3;
  assign xor_cse_482 = Encrypt_Top_sbox_2_and_2_cse_17_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1
      ^ state_4_4_58_lpi_3;
  assign state_4_17_sva_2_mx0w4 = xor_cse_479 ^ xor_cse_480 ^ xor_cse_481 ^ xor_cse_482;
  assign xor_cse_483 = state_2_18_1_lpi_4 ^ (state_4_3_31_0_sva_18 & state_3_3_31_0_sva_18)
      ^ state_4_3_31_0_sva_18 ^ plaintext_31_0_sva_18;
  assign xor_cse_487 = state_4_3_31_0_sva_13 & state_3_3_31_0_sva_13;
  assign xor_cse_488 = state_2_13_1_lpi_4 ^ (state_4_4_13_lpi_3 & state_3_13_lpi_3)
      ^ state_4_4_13_lpi_3 ^ state_1_1_31_0_lpi_4_13;
  assign xor_cse_490 = state_4_4_25_lpi_3 ^ state_1_1_31_0_lpi_4_25 ^ Encrypt_Top_sbox_1_and_cse_25_sva_1
      ^ state_3_25_lpi_3;
  assign xor_cse_491 = state_4_4_18_lpi_3 ^ state_1_1_31_0_lpi_4_18 ^ Encrypt_Top_sbox_1_and_cse_18_sva_1
      ^ state_3_18_lpi_3;
  assign xor_cse_492 = state_1_1_63_32_lpi_4_31 ^ (state_4_4_59_lpi_3 & state_1_1_63_32_lpi_4_31)
      ^ state_3_59_lpi_3 ^ (state_1_1_63_32_lpi_4_31 & state_0_59_lpi_6);
  assign state_4_18_sva_2_mx0w4 = xor_cse_490 ^ xor_cse_491 ^ xor_cse_492 ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1 ^ state_4_4_59_lpi_3;
  assign xor_cse_494 = state_4_3_31_0_sva_14 & state_3_3_31_0_sva_14;
  assign xor_cse_495 = state_4_3_31_0_sva_19 & state_3_3_31_0_sva_19;
  assign xor_cse_496 = state_2_14_1_lpi_4 ^ (state_4_4_14_lpi_3 & state_3_14_lpi_3)
      ^ state_4_4_14_lpi_3 ^ state_1_1_31_0_lpi_4_14;
  assign xor_cse_498 = state_4_4_19_lpi_3 ^ state_1_1_31_0_lpi_4_19 ^ Encrypt_Top_sbox_1_and_cse_19_sva_1
      ^ state_3_19_lpi_3;
  assign xor_cse_499 = state_1_1_63_32_lpi_4_4 ^ (state_4_4_60_lpi_3 & state_1_1_63_32_lpi_4_4)
      ^ state_3_60_lpi_3 ^ (state_1_1_63_32_lpi_4_4 & state_0_60_lpi_6);
  assign xor_cse_500 = state_4_4_26_lpi_3 ^ state_1_1_31_0_lpi_4_26 ^ Encrypt_Top_sbox_1_and_cse_26_sva_1
      ^ state_3_26_lpi_3;
  assign state_4_19_sva_2_mx0w4 = xor_cse_498 ^ xor_cse_499 ^ xor_cse_500 ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_26_sva_1 ^ state_4_4_60_lpi_3;
  assign xor_cse_502 = state_4_3_31_0_sva_15 & state_3_3_31_0_sva_15;
  assign xor_cse_503 = state_4_3_31_0_sva_20 & state_3_3_31_0_sva_20;
  assign xor_cse_504 = state_2_15_1_lpi_4 ^ (state_4_4_15_lpi_3 & state_3_15_lpi_3)
      ^ state_4_4_15_lpi_3 ^ state_1_1_31_0_lpi_4_15;
  assign xor_cse_505 = Encrypt_Top_sbox_1_and_792 ^ state_4_4_20_lpi_3 ^ state_2_20_1_lpi_4
      ^ state_1_1_31_0_lpi_4_20;
  assign xor_cse_506 = state_1_1_63_32_lpi_4_9 ^ (state_4_4_9_lpi_3 & state_1_1_63_32_lpi_4_9)
      ^ state_3_9_lpi_3 ^ (state_1_1_63_32_lpi_4_9 & state_0_9_lpi_6);
  assign xor_cse_507 = state_1_1_63_32_lpi_4_17 ^ state_4_4_43_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_43_sva_1
      ^ state_3_43_lpi_3;
  assign state_4_2_sva_2_mx0w4 = xor_cse_84 ^ xor_cse_506 ^ xor_cse_507 ^ state_4_4_2_lpi_3
      ^ state_4_4_9_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1;
  assign xor_cse_509 = xor_cse_502 ^ state_4_3_31_0_sva_15 ^ state_2_15_1_lpi_4 ^
      plaintext_31_0_sva_15;
  assign xor_cse_511 = state_4_3_31_0_sva_21 & state_3_3_31_0_sva_21;
  assign xor_cse_513 = (state_4_4_21_lpi_3 & state_3_21_lpi_3) ^ state_4_4_21_lpi_3
      ^ state_2_21_1_lpi_4 ^ state_1_1_31_0_lpi_4_21;
  assign xor_cse_514 = state_4_4_20_lpi_3 ^ state_1_1_31_0_lpi_4_20 ^ Encrypt_Top_sbox_1_and_cse_20_sva_1
      ^ state_3_20_lpi_3;
  assign xor_cse_515 = state_1_1_63_32_lpi_4_5 ^ (state_4_4_61_lpi_3 & state_1_1_63_32_lpi_4_5)
      ^ state_3_61_lpi_3 ^ (state_1_1_63_32_lpi_4_5 & state_0_61_lpi_6);
  assign xor_cse_516 = Encrypt_Top_sbox_1_and_cse_27_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_27_sva_1
      ^ state_4_4_27_lpi_3 ^ state_3_27_lpi_3;
  assign state_4_20_sva_2_mx0w4 = xor_cse_514 ^ xor_cse_515 ^ xor_cse_516 ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1
      ^ state_1_1_31_0_lpi_4_27 ^ state_4_4_61_lpi_3;
  assign xor_cse_519 = state_4_3_31_0_sva_22 & state_3_3_31_0_sva_22;
  assign xor_cse_520 = state_4_4_21_lpi_3 ^ state_1_1_31_0_lpi_4_21 ^ Encrypt_Top_sbox_1_and_cse_21_sva_1
      ^ state_3_21_lpi_3;
  assign xor_cse_521 = state_1_1_63_32_lpi_4_6 ^ (state_4_4_62_lpi_3 & state_1_1_63_32_lpi_4_6)
      ^ state_3_62_lpi_3 ^ (state_1_1_63_32_lpi_4_6 & state_0_62_lpi_6);
  assign xor_cse_522 = state_4_4_28_lpi_3 ^ state_1_1_31_0_lpi_4_28 ^ Encrypt_Top_sbox_1_and_cse_28_sva_1
      ^ state_3_28_lpi_3;
  assign state_4_21_sva_2_mx0w4 = xor_cse_520 ^ xor_cse_521 ^ xor_cse_522 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_28_sva_1 ^ state_4_4_62_lpi_3;
  assign xor_cse_525 = state_4_3_31_0_sva_23 & state_3_3_31_0_sva_23;
  assign xor_cse_526 = state_4_4_29_lpi_3 ^ state_1_1_31_0_lpi_4_29 ^ Encrypt_Top_sbox_1_and_cse_29_sva_1
      ^ state_3_29_lpi_3;
  assign xor_cse_527 = state_1_1_63_32_lpi_4_7 ^ (state_4_4_63_lpi_3 & state_1_1_63_32_lpi_4_7)
      ^ state_3_63_lpi_3 ^ (state_1_1_63_32_lpi_4_7 & state_0_63_lpi_6);
  assign xor_cse_528 = state_4_4_22_lpi_3 ^ state_1_1_31_0_lpi_4_22 ^ Encrypt_Top_sbox_1_and_cse_22_sva_1
      ^ state_3_22_lpi_3;
  assign xor_cse_529 = Encrypt_Top_sbox_2_and_2_cse_22_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_29_sva_1
      ^ state_4_4_63_lpi_3;
  assign state_4_22_sva_2_mx0w4 = xor_cse_526 ^ xor_cse_527 ^ xor_cse_528 ^ xor_cse_529;
  assign xor_cse_532 = state_4_3_31_0_sva_24 & state_3_3_31_0_sva_24;
  assign state_4_4_23_sva_1_mx0w4 = xor_cse_56 ^ xor_cse_468 ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_30_sva_1 ^ state_4_4_30_lpi_3 ^ state_3_30_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1 ^ state_1_1_31_0_lpi_4_30 ^ state_4_4_0_lpi_3;
  assign xor_cse_535 = state_4_3_31_0_sva_25 & state_3_3_31_0_sva_25;
  assign xor_cse_536 = state_4_4_31_lpi_3 ^ state_1_1_31_0_lpi_4_31 ^ Encrypt_Top_sbox_1_and_cse_31_sva_1
      ^ state_3_31_lpi_3;
  assign state_4_4_24_sva_1_mx0w4 = xor_cse_70 ^ xor_cse_536 ^ xor_cse_481 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_31_sva_1 ^ state_4_4_1_lpi_3;
  assign xor_cse_538 = state_4_3_31_0_sva_26 & state_3_3_31_0_sva_26;
  assign xor_cse_539 = state_2_26_1_lpi_4 ^ (state_4_4_26_lpi_3 & state_3_26_lpi_3)
      ^ state_4_4_26_lpi_3 ^ state_1_1_31_0_lpi_4_26;
  assign xor_cse_542 = Encrypt_Top_sbox_2_and_2_cse_25_sva_1 ^ state_4_4_32_lpi_3
      ^ state_4_4_2_lpi_3;
  assign state_4_25_sva_2_mx0w4 = xor_cse_84 ^ xor_cse_490 ^ xor_cse_412 ^ xor_cse_542;
  assign xor_cse_543 = state_4_3_31_0_sva_27 & state_3_3_31_0_sva_27;
  assign xor_cse_544 = state_4_4_27_lpi_3 ^ state_1_1_31_0_lpi_4_27 ^ (state_4_4_27_lpi_3
      & state_3_27_lpi_3) ^ state_2_27_1_lpi_4;
  assign xor_cse_546 = Encrypt_Top_sbox_1_and_796 ^ state_4_4_22_lpi_3 ^ state_2_22_1_lpi_4
      ^ state_1_1_31_0_lpi_4_22;
  assign xor_cse_547 = Encrypt_Top_sbox_2_and_2_cse_26_sva_1 ^ state_4_4_33_lpi_3
      ^ state_4_4_3_lpi_3;
  assign state_4_26_sva_2_mx0w4 = xor_cse_102 ^ xor_cse_425 ^ xor_cse_500 ^ xor_cse_547;
  assign xor_cse_548 = state_4_3_31_0_sva_28 & state_3_3_31_0_sva_28;
  assign xor_cse_549 = state_2_28_1_lpi_4 ^ state_4_4_28_lpi_3 ^ state_1_1_31_0_lpi_4_28
      ^ Encrypt_Top_sbox_1_and_808;
  assign xor_cse_551 = Encrypt_Top_sbox_1_and_798 ^ state_4_4_23_lpi_3 ^ state_2_23_1_lpi_4
      ^ state_1_1_31_0_lpi_4_23;
  assign xor_cse_552 = state_1_1_31_0_lpi_4_27 ^ state_4_4_34_lpi_3 ^ state_4_4_4_lpi_3;
  assign state_4_27_sva_2_mx0w4 = xor_cse_111 ^ xor_cse_439 ^ xor_cse_516 ^ xor_cse_552;
  assign xor_cse_553 = state_4_3_31_0_sva_29 & state_3_3_31_0_sva_29;
  assign xor_cse_554 = state_2_29_1_lpi_4 ^ (state_4_4_29_lpi_3 & state_3_29_lpi_3)
      ^ state_4_4_29_lpi_3 ^ state_1_1_31_0_lpi_4_29;
  assign xor_cse_556 = Encrypt_Top_sbox_1_and_800 ^ state_4_4_24_lpi_3 ^ state_2_24_1_lpi_4
      ^ state_1_1_31_0_lpi_4_24;
  assign xor_cse_557 = Encrypt_Top_sbox_2_and_2_cse_28_sva_1 ^ state_4_4_35_lpi_3
      ^ state_4_4_5_lpi_3;
  assign state_4_28_sva_2_mx0w4 = xor_cse_124 ^ xor_cse_458 ^ xor_cse_522 ^ xor_cse_557;
  assign xor_cse_558 = state_4_3_31_0_sva_30 & state_3_3_31_0_sva_30;
  assign xor_cse_559 = state_4_4_30_lpi_3 ^ state_1_1_31_0_lpi_4_30 ^ (state_4_4_30_lpi_3
      & state_3_30_lpi_3) ^ state_2_30_1_lpi_4;
  assign xor_cse_561 = Encrypt_Top_sbox_1_and_802 ^ state_4_4_25_lpi_3 ^ state_2_25_1_lpi_4
      ^ state_1_1_31_0_lpi_4_25;
  assign xor_cse_562 = xor_cse_136 ^ state_4_4_6_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_29_sva_1
      ^ state_4_4_36_lpi_3;
  assign state_4_29_sva_2_mx0w4 = xor_cse_562 ^ xor_cse_526 ^ Encrypt_Top_sbox_3_and_cse_36_sva_1
      ^ state_3_36_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1 ^ state_1_1_63_32_lpi_4_10;
  assign xor_cse_565 = state_4_3_31_0_sva_31 & state_3_3_31_0_sva_31;
  assign xor_cse_566 = state_2_31_1_lpi_4 ^ (state_4_4_31_lpi_3 & state_3_31_lpi_3)
      ^ state_4_4_31_lpi_3 ^ state_1_1_31_0_lpi_4_31;
  assign xor_cse_568 = state_1_1_63_32_lpi_4_18 ^ (state_4_4_44_lpi_3 & state_1_1_63_32_lpi_4_18)
      ^ state_3_44_lpi_3 ^ (state_1_1_63_32_lpi_4_18 & state_0_44_lpi_6);
  assign xor_cse_569 = Encrypt_Top_sbox_1_and_cse_10_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_10_sva_1
      ^ state_4_4_10_lpi_3 ^ state_3_10_lpi_3;
  assign xor_cse_570 = xor_cse_102 ^ state_4_4_3_lpi_3 ^ state_1_1_31_0_lpi_4_10
      ^ state_4_4_44_lpi_3;
  assign state_4_3_sva_2_mx0w4 = xor_cse_568 ^ xor_cse_569 ^ xor_cse_570;
  assign xor_cse_571 = state_4_3_63_32_sva_0 ^ (state_4_3_63_32_sva_0 & state_3_3_63_32_sva_0)
      ^ state_2_32_1_lpi_4 ^ plaintext_63_32_sva_0;
  assign xor_cse_574 = xor_cse_543 ^ state_4_3_31_0_sva_27 ^ state_2_27_1_lpi_4 ^
      plaintext_31_0_sva_27;
  assign xor_cse_575 = state_2_32_1_lpi_4 ^ Encrypt_Top_sbox_1_and_816 ^ state_4_4_32_lpi_3
      ^ state_1_1_63_32_lpi_4_0;
  assign xor_cse_576 = Encrypt_Top_sbox_1_and_816 ^ state_4_4_32_lpi_3 ^ state_2_32_1_lpi_4
      ^ state_1_1_31_0_lpi_4_8;
  assign xor_cse_577 = xor_cse_148 ^ state_4_4_7_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_30_sva_1
      ^ state_4_4_30_lpi_3;
  assign state_4_30_sva_2_mx0w5 = xor_cse_577 ^ state_3_30_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1
      ^ state_1_1_31_0_lpi_4_30 ^ Encrypt_Top_sbox_3_and_cse_37_sva_1 ^ state_4_4_37_lpi_3
      ^ state_3_37_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1 ^ state_1_1_63_32_lpi_4_11;
  assign xor_cse_581 = state_2_33_1_lpi_4 ^ plaintext_63_32_sva_1 ^ (state_4_3_63_32_sva_1
      & state_3_3_63_32_sva_1) ^ state_4_3_63_32_sva_1;
  assign xor_cse_585 = state_2_33_1_lpi_4 ^ Encrypt_Top_sbox_1_and_818 ^ state_4_4_33_lpi_3
      ^ state_1_1_63_32_lpi_4_1;
  assign xor_cse_586 = state_4_4_33_lpi_3 ^ Encrypt_Top_sbox_1_and_818 ^ state_2_33_1_lpi_4
      ^ state_1_1_31_0_lpi_4_9;
  assign xor_cse_587 = state_1_1_63_32_lpi_4_8 ^ (state_4_4_8_lpi_3 & state_1_1_63_32_lpi_4_8)
      ^ state_3_8_lpi_3 ^ (state_1_1_63_32_lpi_4_8 & state_0_8_lpi_6);
  assign xor_cse_588 = state_1_1_63_32_lpi_4_12 ^ (state_4_4_38_lpi_3 & state_1_1_63_32_lpi_4_12)
      ^ state_3_38_lpi_3 ^ (state_1_1_63_32_lpi_4_12 & state_0_38_lpi_6);
  assign xor_cse_589 = Encrypt_Top_sbox_2_and_2_cse_31_sva_1 ^ state_4_4_38_lpi_3
      ^ state_4_4_8_lpi_3;
  assign state_4_31_sva_2_mx0w5 = xor_cse_536 ^ xor_cse_587 ^ xor_cse_588 ^ xor_cse_589;
  assign xor_cse_590 = state_4_3_63_32_sva_2 & state_3_3_63_32_sva_2;
  assign xor_cse_591 = state_2_34_1_lpi_4 ^ Encrypt_Top_sbox_1_and_820 ^ state_4_4_34_lpi_3
      ^ Encrypt_Top_sbox_1_and_808;
  assign xor_cse_594 = state_4_4_11_lpi_3 ^ state_1_1_31_0_lpi_4_11 ^ Encrypt_Top_sbox_1_and_cse_11_sva_1
      ^ state_3_11_lpi_3;
  assign xor_cse_595 = state_1_1_63_32_lpi_4_19 ^ Encrypt_Top_sbox_3_and_cse_45_sva_1
      ^ state_4_4_45_lpi_3 ^ state_3_45_lpi_3;
  assign state_4_4_sva_2_mx0w5 = xor_cse_111 ^ xor_cse_594 ^ xor_cse_595 ^ state_4_4_4_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1;
  assign xor_cse_597 = state_4_3_63_32_sva_3 ^ (state_4_3_63_32_sva_3 & state_3_3_63_32_sva_3)
      ^ state_2_35_1_lpi_4 ^ plaintext_63_32_sva_3;
  assign xor_cse_601 = state_2_35_1_lpi_4 ^ Encrypt_Top_sbox_1_and_822 ^ state_4_4_35_lpi_3
      ^ state_1_1_63_32_lpi_4_3;
  assign xor_cse_602 = state_4_4_35_lpi_3 ^ Encrypt_Top_sbox_1_and_822 ^ state_2_35_1_lpi_4
      ^ state_1_1_63_32_lpi_4_1;
  assign xor_cse_603 = state_4_4_12_lpi_3 ^ state_1_1_31_0_lpi_4_12 ^ Encrypt_Top_sbox_1_and_cse_12_sva_1
      ^ state_3_12_lpi_3;
  assign xor_cse_604 = state_1_1_63_32_lpi_4_2 ^ (state_4_4_46_lpi_3 & state_1_1_63_32_lpi_4_2)
      ^ state_3_46_lpi_3 ^ (state_1_1_63_32_lpi_4_2 & state_0_46_lpi_6);
  assign xor_cse_605 = state_4_4_5_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_12_sva_1
      ^ state_4_4_46_lpi_3;
  assign state_4_5_sva_2_mx0w5 = xor_cse_124 ^ xor_cse_603 ^ xor_cse_604 ^ xor_cse_605;
  assign xor_cse_606 = state_4_3_63_32_sva_4 & state_3_3_63_32_sva_4;
  assign xor_cse_607 = Encrypt_Top_sbox_1_and_824 ^ state_4_4_36_lpi_3 ^ state_2_36_1_lpi_4
      ^ state_1_1_63_32_lpi_4_4;
  assign xor_cse_608 = state_1_1_63_32_lpi_4_10 ^ state_4_4_36_lpi_3 ^ Encrypt_Top_sbox_1_and_824
      ^ state_2_36_1_lpi_4;
  assign xor_cse_609 = state_4_4_13_lpi_3 ^ state_1_1_31_0_lpi_4_13 ^ Encrypt_Top_sbox_1_and_cse_13_sva_1
      ^ state_3_13_lpi_3;
  assign xor_cse_610 = state_1_1_63_32_lpi_4_20 ^ Encrypt_Top_sbox_3_and_cse_47_sva_1
      ^ state_4_4_47_lpi_3 ^ state_3_47_lpi_3;
  assign state_4_6_sva_2_mx0w5 = xor_cse_136 ^ xor_cse_609 ^ xor_cse_610 ^ state_4_4_6_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1;
  assign xor_cse_614 = state_4_3_63_32_sva_5 & state_3_3_63_32_sva_5;
  assign xor_cse_613 = xor_cse_614 ^ state_4_3_63_32_sva_5 ^ state_2_37_1_lpi_4 ^
      plaintext_63_32_sva_5;
  assign xor_cse_616 = state_1_1_63_32_lpi_4_11 ^ state_4_4_37_lpi_3 ^ Encrypt_Top_sbox_1_and_826
      ^ state_2_37_1_lpi_4;
  assign xor_cse_618 = state_4_4_14_lpi_3 ^ state_1_1_31_0_lpi_4_14 ^ Encrypt_Top_sbox_1_and_cse_14_sva_1
      ^ state_3_14_lpi_3;
  assign xor_cse_619 = state_1_1_63_32_lpi_4_21 ^ Encrypt_Top_sbox_3_and_cse_48_sva_1
      ^ state_4_4_48_lpi_3 ^ state_3_48_lpi_3;
  assign state_4_7_sva_2_mx0w5 = xor_cse_148 ^ xor_cse_618 ^ xor_cse_619 ^ state_4_4_7_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1;
  assign xor_cse_621 = state_4_3_63_32_sva_6 ^ (state_4_3_63_32_sva_6 & state_3_3_63_32_sva_6)
      ^ state_2_38_1_lpi_4 ^ plaintext_63_32_sva_6;
  assign xor_cse_624 = state_1_1_63_32_lpi_4_12 ^ state_2_38_1_lpi_4 ^ Encrypt_Top_sbox_1_and_828
      ^ state_4_4_38_lpi_3;
  assign state_4_32_sva_2_mx0w5 = xor_cse_412 ^ xor_cse_506 ^ state_4_4_32_lpi_3
      ^ Encrypt_Top_sbox_3_and_cse_39_sva_1 ^ state_4_4_39_lpi_3 ^ state_3_39_lpi_3
      ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1 ^ state_1_1_63_32_lpi_4_13 ^ state_4_4_9_lpi_3;
  assign xor_cse_628 = xor_cse_590 ^ state_4_3_63_32_sva_2 ^ state_2_34_1_lpi_4 ^
      plaintext_63_32_sva_2;
  assign xor_cse_629 = (state_4_3_63_32_sva_7 & state_3_3_63_32_sva_7) ^ state_4_3_63_32_sva_7
      ^ state_2_39_1_lpi_4 ^ plaintext_63_32_sva_7;
  assign xor_cse_631 = state_4_4_34_lpi_3 ^ Encrypt_Top_sbox_1_and_820 ^ state_2_34_1_lpi_4
      ^ state_1_1_63_32_lpi_4_2;
  assign xor_cse_633 = state_1_1_63_32_lpi_4_13 ^ state_4_4_39_lpi_3 ^ Encrypt_Top_sbox_1_and_830
      ^ state_2_39_1_lpi_4;
  assign xor_cse_634 = Encrypt_Top_sbox_1_and_820 ^ state_4_4_34_lpi_3 ^ state_2_34_1_lpi_4
      ^ state_1_1_63_32_lpi_4_0;
  assign xor_cse_635 = state_1_1_63_32_lpi_4_14 ^ (state_4_4_40_lpi_3 & state_1_1_63_32_lpi_4_14)
      ^ state_3_40_lpi_3 ^ (state_1_1_63_32_lpi_4_14 & state_0_40_lpi_6);
  assign xor_cse_636 = state_4_4_33_lpi_3 ^ state_4_4_40_lpi_3 ^ state_1_1_31_0_lpi_4_10;
  assign state_4_33_sva_2_mx0w5 = xor_cse_425 ^ xor_cse_635 ^ xor_cse_569 ^ xor_cse_636;
  assign xor_cse_637 = state_4_3_63_32_sva_8 ^ (state_4_3_63_32_sva_8 & state_3_3_63_32_sva_8)
      ^ state_2_40_1_lpi_4 ^ plaintext_63_32_sva_8;
  assign xor_cse_641 = state_1_1_63_32_lpi_4_14 ^ state_2_40_1_lpi_4 ^ Encrypt_Top_sbox_1_and_832
      ^ state_4_4_40_lpi_3;
  assign xor_cse_643 = state_4_4_41_lpi_3 ^ state_3_41_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_41_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_41_sva_1;
  assign state_4_34_sva_2_mx0w5 = xor_cse_594 ^ xor_cse_439 ^ xor_cse_643 ^ state_4_4_34_lpi_3
      ^ state_1_1_63_32_lpi_4_15 ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1;
  assign xor_cse_645 = state_4_3_63_32_sva_9 ^ (state_4_3_63_32_sva_9 & state_3_3_63_32_sva_9)
      ^ state_2_41_1_lpi_4 ^ plaintext_63_32_sva_9;
  assign xor_cse_650 = state_1_1_63_32_lpi_4_15 ^ state_4_4_41_lpi_3 ^ Encrypt_Top_sbox_1_and_834
      ^ state_2_41_1_lpi_4;
  assign xor_cse_651 = state_1_1_63_32_lpi_4_16 ^ (state_4_4_42_lpi_3 & state_1_1_63_32_lpi_4_16)
      ^ state_3_42_lpi_3 ^ (state_1_1_63_32_lpi_4_16 & state_0_42_lpi_6);
  assign state_4_35_sva_2_mx0w5 = xor_cse_603 ^ xor_cse_651 ^ xor_cse_458 ^ state_4_4_35_lpi_3
      ^ state_4_4_42_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_12_sva_1;
  assign xor_cse_653 = state_4_3_63_32_sva_10 & state_3_3_63_32_sva_10;
  assign xor_cse_656 = state_1_1_63_32_lpi_4_16 ^ state_2_42_1_lpi_4 ^ Encrypt_Top_sbox_1_and_836
      ^ state_4_4_42_lpi_3;
  assign state_4_36_sva_2_mx0w5 = xor_cse_609 ^ xor_cse_507 ^ Encrypt_Top_sbox_3_and_cse_36_sva_1
      ^ state_4_4_36_lpi_3 ^ state_3_36_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1
      ^ state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1;
  assign xor_cse_659 = state_4_3_63_32_sva_11 ^ (state_4_3_63_32_sva_11 & state_3_3_63_32_sva_11)
      ^ state_2_43_1_lpi_4 ^ plaintext_63_32_sva_11;
  assign xor_cse_664 = state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_1_and_838 ^ state_4_4_43_lpi_3
      ^ state_2_43_1_lpi_4;
  assign state_4_37_sva_2_mx0w5 = xor_cse_618 ^ xor_cse_568 ^ Encrypt_Top_sbox_3_and_cse_37_sva_1
      ^ state_4_4_37_lpi_3 ^ state_3_37_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1
      ^ state_1_1_63_32_lpi_4_11 ^ state_4_4_44_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1;
  assign xor_cse_667 = state_4_3_63_32_sva_12 ^ (state_4_3_63_32_sva_12 & state_3_3_63_32_sva_12)
      ^ state_2_44_1_lpi_4 ^ plaintext_63_32_sva_12;
  assign xor_cse_672 = state_1_1_63_32_lpi_4_18 ^ state_2_44_1_lpi_4 ^ Encrypt_Top_sbox_1_and_840
      ^ state_4_4_44_lpi_3;
  assign xor_cse_673 = state_4_4_15_lpi_3 ^ state_1_1_31_0_lpi_4_15 ^ Encrypt_Top_sbox_1_and_cse_15_sva_1
      ^ state_3_15_lpi_3;
  assign state_4_38_sva_2_mx0w5 = xor_cse_673 ^ xor_cse_588 ^ xor_cse_595 ^ state_4_4_38_lpi_3
      ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1;
  assign xor_cse_676 = (state_4_3_63_32_sva_13 & state_3_3_63_32_sva_13) ^ state_4_3_63_32_sva_13
      ^ state_2_45_1_lpi_4 ^ plaintext_63_32_sva_13;
  assign xor_cse_680 = state_1_1_63_32_lpi_4_19 ^ state_4_4_45_lpi_3 ^ Encrypt_Top_sbox_1_and_842
      ^ state_2_45_1_lpi_4;
  assign state_4_39_sva_2_mx0w5 = xor_cse_469 ^ xor_cse_604 ^ Encrypt_Top_sbox_3_and_cse_39_sva_1
      ^ state_4_4_39_lpi_3 ^ state_3_39_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1
      ^ state_1_1_63_32_lpi_4_13 ^ state_4_4_46_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1;
  assign xor_cse_683 = state_4_3_63_32_sva_14 ^ (state_4_3_63_32_sva_14 & state_3_3_63_32_sva_14)
      ^ state_2_46_1_lpi_4 ^ plaintext_63_32_sva_14;
  assign xor_cse_685 = state_4_4_46_lpi_3 ^ Encrypt_Top_sbox_1_and_844 ^ state_2_46_1_lpi_4
      ^ xor_cse_641;
  assign state_4_40_sva_2_mx0w5 = xor_cse_479 ^ xor_cse_635 ^ xor_cse_610 ^ state_4_4_40_lpi_3
      ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_17_sva_1;
  assign xor_cse_689 = xor_cse_653 ^ state_4_3_63_32_sva_10 ^ state_2_42_1_lpi_4
      ^ plaintext_63_32_sva_10;
  assign xor_cse_691 = state_4_3_63_32_sva_15 & state_3_3_63_32_sva_15;
  assign xor_cse_690 = xor_cse_691 ^ state_4_3_63_32_sva_15 ^ state_2_47_1_lpi_4
      ^ plaintext_63_32_sva_15;
  assign xor_cse_694 = state_1_1_63_32_lpi_4_20 ^ state_4_4_47_lpi_3 ^ Encrypt_Top_sbox_1_and_846
      ^ state_2_47_1_lpi_4;
  assign state_4_41_sva_2_mx0w5 = xor_cse_491 ^ xor_cse_643 ^ xor_cse_619 ^ state_1_1_63_32_lpi_4_15
      ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1;
  assign xor_cse_698 = state_4_3_63_32_sva_16 & state_3_3_63_32_sva_16;
  assign xor_cse_701 = state_1_1_63_32_lpi_4_21 ^ state_4_4_48_lpi_3 ^ Encrypt_Top_sbox_1_and_848
      ^ state_2_48_1_lpi_4;
  assign xor_cse_702 = state_1_1_63_32_lpi_4_22 ^ (state_4_4_49_lpi_3 & state_1_1_63_32_lpi_4_22)
      ^ state_3_49_lpi_3 ^ (state_1_1_63_32_lpi_4_22 & state_0_49_lpi_6);
  assign state_4_42_sva_2_mx0w5 = xor_cse_498 ^ xor_cse_651 ^ xor_cse_702 ^ state_4_4_42_lpi_3
      ^ state_4_4_49_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1;
  assign xor_cse_705 = state_4_3_63_32_sva_17 & state_3_3_63_32_sva_17;
  assign xor_cse_708 = state_1_1_63_32_lpi_4_22 ^ state_2_49_1_lpi_4 ^ Encrypt_Top_sbox_1_and_850
      ^ state_4_4_49_lpi_3;
  assign xor_cse_709 = state_4_4_50_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_50_sva_1 ^
      state_3_50_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_50_sva_1;
  assign state_4_43_sva_2_mx0w5 = xor_cse_514 ^ xor_cse_507 ^ xor_cse_709 ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1
      ^ state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1;
  assign xor_cse_713 = state_4_3_63_32_sva_18 & state_3_3_63_32_sva_18;
  assign xor_cse_716 = state_1_1_63_32_lpi_4_23 ^ state_4_4_50_lpi_3 ^ Encrypt_Top_sbox_1_and_852
      ^ state_2_50_1_lpi_4;
  assign xor_cse_717 = state_1_1_63_32_lpi_4_24 ^ (state_4_4_51_lpi_3 & state_1_1_63_32_lpi_4_24)
      ^ state_3_51_lpi_3 ^ (state_1_1_63_32_lpi_4_24 & state_0_51_lpi_6);
  assign state_4_44_sva_2_mx0w5 = xor_cse_520 ^ xor_cse_568 ^ xor_cse_717 ^ state_4_4_44_lpi_3
      ^ state_4_4_51_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1;
  assign xor_cse_721 = state_4_3_63_32_sva_19 & state_3_3_63_32_sva_19;
  assign xor_cse_722 = state_2_46_1_lpi_4 ^ Encrypt_Top_sbox_1_and_844 ^ state_4_4_46_lpi_3
      ^ state_1_1_63_32_lpi_4_14;
  assign xor_cse_724 = state_1_1_63_32_lpi_4_24 ^ state_2_51_1_lpi_4 ^ Encrypt_Top_sbox_1_and_854
      ^ state_4_4_51_lpi_3;
  assign xor_cse_725 = Encrypt_Top_sbox_1_and_844 ^ state_4_4_46_lpi_3 ^ state_2_46_1_lpi_4
      ^ state_1_1_63_32_lpi_4_2;
  assign xor_cse_726 = state_1_1_63_32_lpi_4_25 ^ (state_4_4_52_lpi_3 & state_1_1_63_32_lpi_4_25)
      ^ state_3_52_lpi_3 ^ (state_1_1_63_32_lpi_4_25 & state_0_52_lpi_6);
  assign state_4_45_sva_2_mx0w5 = xor_cse_528 ^ xor_cse_726 ^ xor_cse_595 ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1
      ^ state_4_4_52_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_22_sva_1;
  assign xor_cse_730 = state_4_3_63_32_sva_20 & state_3_3_63_32_sva_20;
  assign xor_cse_732 = state_1_1_63_32_lpi_4_25 ^ state_2_52_1_lpi_4 ^ Encrypt_Top_sbox_1_and_856
      ^ state_4_4_52_lpi_3;
  assign xor_cse_734 = state_1_1_63_32_lpi_4_26 ^ (state_4_4_53_lpi_3 & state_1_1_63_32_lpi_4_26)
      ^ state_3_53_lpi_3 ^ (state_1_1_63_32_lpi_4_26 & state_0_53_lpi_6);
  assign xor_cse_735 = state_4_4_46_lpi_3 ^ state_4_4_53_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1;
  assign state_4_46_sva_2_mx0w5 = xor_cse_468 ^ xor_cse_604 ^ xor_cse_734 ^ xor_cse_735;
  assign xor_cse_736 = state_4_3_63_32_sva_21 & state_3_3_63_32_sva_21;
  assign xor_cse_739 = state_1_1_63_32_lpi_4_26 ^ state_2_53_1_lpi_4 ^ Encrypt_Top_sbox_1_and_858
      ^ state_4_4_53_lpi_3;
  assign xor_cse_740 = state_1_1_63_32_lpi_4_27 ^ (state_4_4_54_lpi_3 & state_1_1_63_32_lpi_4_27)
      ^ state_3_54_lpi_3 ^ (state_1_1_63_32_lpi_4_27 & state_0_54_lpi_6);
  assign state_4_47_sva_2_mx0w5 = xor_cse_740 ^ xor_cse_481 ^ xor_cse_610 ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1
      ^ state_4_4_54_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1;
  assign xor_cse_742 = state_4_3_63_32_sva_22 & state_3_3_63_32_sva_22;
  assign xor_cse_743 = state_4_4_54_lpi_3 ^ Encrypt_Top_sbox_1_and_860 ^ state_2_54_1_lpi_4
      ^ xor_cse_708;
  assign xor_cse_746 = state_1_1_63_32_lpi_4_28 ^ (state_4_4_55_lpi_3 & state_1_1_63_32_lpi_4_28)
      ^ state_3_55_lpi_3 ^ (state_1_1_63_32_lpi_4_28 & state_0_55_lpi_6);
  assign state_4_48_sva_2_mx0w5 = xor_cse_490 ^ xor_cse_746 ^ xor_cse_619 ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1
      ^ state_4_4_55_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1;
  assign xor_cse_748 = state_4_3_63_32_sva_23 & state_3_3_63_32_sva_23;
  assign xor_cse_749 = state_2_55_1_lpi_4 ^ Encrypt_Top_sbox_1_and_862 ^ state_4_4_55_lpi_3
      ^ xor_cse_716;
  assign xor_cse_752 = state_1_1_63_32_lpi_4_29 ^ (state_4_4_56_lpi_3 & state_1_1_63_32_lpi_4_29)
      ^ state_3_56_lpi_3 ^ (state_1_1_63_32_lpi_4_29 & state_0_56_lpi_6);
  assign xor_cse_753 = state_4_4_49_lpi_3 ^ state_4_4_56_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_26_sva_1;
  assign state_4_49_sva_2_mx0w5 = xor_cse_752 ^ xor_cse_702 ^ xor_cse_500 ^ xor_cse_753;
  assign xor_cse_754 = state_4_3_63_32_sva_24 & state_3_3_63_32_sva_24;
  assign xor_cse_755 = state_4_4_56_lpi_3 ^ state_2_56_1_lpi_4 ^ Encrypt_Top_sbox_1_and_864
      ^ xor_cse_724;
  assign state_4_50_sva_2_mx0w5 = xor_cse_470 ^ xor_cse_516 ^ xor_cse_709 ^ state_1_1_63_32_lpi_4_23
      ^ state_4_4_57_lpi_3 ^ state_1_1_31_0_lpi_4_27;
  assign xor_cse_759 = state_4_3_63_32_sva_25 & state_3_3_63_32_sva_25;
  assign xor_cse_760 = state_2_57_1_lpi_4 ^ state_4_4_57_lpi_3 ^ Encrypt_Top_sbox_1_and_866
      ^ xor_cse_732;
  assign xor_cse_763 = state_4_4_51_lpi_3 ^ state_4_4_58_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_28_sva_1;
  assign state_4_51_sva_2_mx0w5 = xor_cse_480 ^ xor_cse_522 ^ xor_cse_717 ^ xor_cse_763;
  assign xor_cse_764 = state_4_3_63_32_sva_26 & state_3_3_63_32_sva_26;
  assign xor_cse_767 = state_2_58_1_lpi_4 ^ Encrypt_Top_sbox_1_and_868 ^ state_4_4_58_lpi_3
      ^ state_1_1_63_32_lpi_4_30;
  assign state_4_52_sva_2_mx0w5 = xor_cse_526 ^ xor_cse_492 ^ xor_cse_726 ^ state_4_4_52_lpi_3
      ^ state_4_4_59_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_29_sva_1;
  assign xor_cse_769 = state_4_3_63_32_sva_27 & state_3_3_63_32_sva_27;
  assign xor_cse_770 = state_1_1_63_32_lpi_4_27 ^ state_4_4_59_lpi_3 ^ Encrypt_Top_sbox_1_and_870
      ^ state_2_59_1_lpi_4;
  assign xor_cse_771 = state_2_54_1_lpi_4 ^ Encrypt_Top_sbox_1_and_860 ^ state_4_4_54_lpi_3
      ^ state_1_1_63_32_lpi_4_22;
  assign xor_cse_775 = state_3_30_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1 ^
      state_1_1_31_0_lpi_4_30;
  assign state_4_53_sva_2_mx0w5 = xor_cse_499 ^ xor_cse_734 ^ state_4_4_53_lpi_3
      ^ state_4_4_60_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_30_sva_1 ^ state_4_4_30_lpi_3
      ^ xor_cse_775;
  assign xor_cse_776 = state_4_3_63_32_sva_28 & state_3_3_63_32_sva_28;
  assign xor_cse_777 = state_1_1_63_32_lpi_4_28 ^ state_4_4_60_lpi_3 ^ Encrypt_Top_sbox_1_and_872
      ^ state_2_60_1_lpi_4;
  assign state_4_54_sva_2_mx0w5 = xor_cse_536 ^ xor_cse_740 ^ xor_cse_515 ^ state_4_4_54_lpi_3
      ^ state_4_4_61_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_31_sva_1;
  assign xor_cse_782 = state_4_3_63_32_sva_29 & state_3_3_63_32_sva_29;
  assign xor_cse_783 = state_1_1_63_32_lpi_4_29 ^ state_4_4_61_lpi_3 ^ Encrypt_Top_sbox_1_and_874
      ^ state_2_61_1_lpi_4;
  assign xor_cse_784 = state_2_55_1_lpi_4 ^ Encrypt_Top_sbox_1_and_862 ^ state_4_4_55_lpi_3
      ^ Encrypt_Top_sbox_1_and_864;
  assign state_4_55_sva_2_mx0w5 = xor_cse_412 ^ xor_cse_746 ^ xor_cse_521 ^ state_4_4_55_lpi_3
      ^ state_4_4_62_lpi_3 ^ state_4_4_32_lpi_3;
  assign xor_cse_788 = state_4_3_63_32_sva_30 & state_3_3_63_32_sva_30;
  assign xor_cse_789 = state_1_1_63_32_lpi_4_30 ^ state_4_4_62_lpi_3 ^ Encrypt_Top_sbox_1_and_876
      ^ state_2_62_1_lpi_4;
  assign xor_cse_790 = state_2_56_1_lpi_4 ^ Encrypt_Top_sbox_1_and_864 ^ state_4_4_56_lpi_3
      ^ Encrypt_Top_sbox_1_and_866;
  assign xor_cse_792 = state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_1_and_876 ^ state_4_4_62_lpi_3
      ^ state_2_62_1_lpi_4;
  assign xor_cse_794 = state_4_4_56_lpi_3 ^ state_4_4_63_lpi_3 ^ state_4_4_33_lpi_3;
  assign state_4_56_sva_2_mx0w5 = xor_cse_425 ^ xor_cse_527 ^ xor_cse_752 ^ xor_cse_794;
  assign xor_cse_795 = state_4_3_63_32_sva_31 & state_3_3_63_32_sva_31;
  assign xor_cse_796 = state_1_1_63_32_lpi_4_31 ^ Encrypt_Top_sbox_1_and_878 ^ state_4_4_63_lpi_3
      ^ state_2_63_1_lpi_4;
  assign xor_cse_797 = state_2_58_1_lpi_4 ^ Encrypt_Top_sbox_1_and_868 ^ state_4_4_58_lpi_3
      ^ state_1_1_63_32_lpi_4_26;
  assign xor_cse_799 = state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_1_and_878 ^ state_4_4_63_lpi_3
      ^ state_2_63_1_lpi_4;
  assign xor_cse_801 = state_4_4_57_lpi_3 ^ state_4_4_0_lpi_3 ^ state_4_4_34_lpi_3;
  assign state_4_57_sva_2_mx0w5 = xor_cse_56 ^ xor_cse_470 ^ xor_cse_439 ^ xor_cse_801;
  assign xor_cse_802 = state_2_0_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0])
      ^ (state_4_3_31_0_sva_0 & state_3_3_31_0_sva_0) ^ state_4_3_31_0_sva_0;
  assign xor_cse_805 = xor_cse_769 ^ state_4_3_63_32_sva_27 ^ state_2_59_1_lpi_4
      ^ plaintext_63_32_sva_27;
  assign xor_cse_806 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]) ^ Encrypt_Top_sbox_1_and_756
      ^ state_4_4_0_lpi_3 ^ state_1_1_31_0_lpi_4_0;
  assign xor_cse_807 = Encrypt_Top_sbox_1_and_870 ^ state_4_4_59_lpi_3 ^ state_2_59_1_lpi_4
      ^ state_1_1_63_32_lpi_4_31;
  assign xor_cse_808 = Encrypt_Top_sbox_1_and_756 ^ state_4_4_0_lpi_3 ^ state_2_0_1_lpi_4
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0]);
  assign xor_cse_809 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1])
      ^ (state_4_3_31_0_sva_1 & state_3_3_31_0_sva_1) ^ state_4_3_31_0_sva_1;
  assign xor_cse_812 = xor_cse_776 ^ state_4_3_63_32_sva_28 ^ state_2_60_1_lpi_4
      ^ plaintext_63_32_sva_28;
  assign xor_cse_813 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]) ^ Encrypt_Top_sbox_1_and_758
      ^ state_4_4_1_lpi_3 ^ state_1_1_31_0_lpi_4_1;
  assign xor_cse_814 = state_2_1_1_lpi_4 ^ Encrypt_Top_sbox_1_and_758 ^ state_4_4_1_lpi_3
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1]);
  assign xor_cse_817 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ (state_4_3_31_0_sva_2 & state_3_3_31_0_sva_2) ^ state_4_3_31_0_sva_2;
  assign xor_cse_820 = xor_cse_782 ^ state_4_3_63_32_sva_29 ^ state_2_61_1_lpi_4
      ^ plaintext_63_32_sva_29;
  assign xor_cse_821 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]) ^ Encrypt_Top_sbox_1_and_760
      ^ state_4_4_2_lpi_3 ^ state_1_1_31_0_lpi_4_2;
  assign xor_cse_822 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ (state_4_3_31_0_sva_3 & state_3_3_31_0_sva_3) ^ state_4_3_31_0_sva_3;
  assign xor_cse_825 = xor_cse_788 ^ state_4_3_63_32_sva_30 ^ state_2_62_1_lpi_4
      ^ plaintext_63_32_sva_30;
  assign xor_cse_826 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]) ^ Encrypt_Top_sbox_1_and_762
      ^ state_4_4_3_lpi_3 ^ state_1_1_31_0_lpi_4_3;
  assign xor_cse_827 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ Encrypt_Top_sbox_1_and_762 ^ state_4_4_3_lpi_3;
  assign xor_cse_829 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4])
      ^ (state_4_3_31_0_sva_4 & state_3_3_31_0_sva_4) ^ state_4_3_31_0_sva_4;
  assign xor_cse_832 = xor_cse_795 ^ state_4_3_63_32_sva_31 ^ state_2_63_1_lpi_4
      ^ plaintext_63_32_sva_31;
  assign xor_cse_833 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]) ^ Encrypt_Top_sbox_1_and_764
      ^ state_4_4_4_lpi_3 ^ state_1_1_31_0_lpi_4_4;
  assign xor_cse_834 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4])
      ^ Encrypt_Top_sbox_1_and_764 ^ state_4_4_4_lpi_3;
  assign xor_cse_835 = state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5])
      ^ (state_4_3_31_0_sva_5 & state_3_3_31_0_sva_5) ^ state_4_3_31_0_sva_5;
  assign xor_cse_839 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]) ^ Encrypt_Top_sbox_1_and_766
      ^ state_4_4_5_lpi_3 ^ state_1_1_31_0_lpi_4_5;
  assign xor_cse_842 = state_2_5_1_lpi_4 ^ Encrypt_Top_sbox_1_and_766 ^ state_4_4_5_lpi_3
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5]);
  assign xor_cse_845 = state_4_3_31_0_sva_8 ^ (state_4_3_31_0_sva_8 & state_3_3_31_0_sva_8)
      ^ state_2_8_1_lpi_4 ^ plaintext_31_0_sva_8;
  assign xor_cse_847 = state_4_3_31_0_sva_9 ^ (state_4_3_31_0_sva_9 & state_3_3_31_0_sva_9)
      ^ state_2_9_1_lpi_4 ^ plaintext_31_0_sva_9;
  assign xor_cse_850 = state_2_8_1_lpi_4 ^ Encrypt_Top_sbox_1_and_880 ^ state_4_4_8_lpi_3
      ^ state_1_1_31_0_lpi_4_8;
  assign xor_cse_851 = state_1_1_31_0_lpi_4_9 ^ Encrypt_Top_sbox_1_and_882 ^ state_4_4_9_lpi_3
      ^ state_2_9_1_lpi_4;
  assign xor_cse_852 = state_2_9_1_lpi_4 ^ Encrypt_Top_sbox_1_and_882 ^ state_4_4_9_lpi_3
      ^ state_1_1_63_32_lpi_4_9;
  assign xor_cse_854 = state_4_4_8_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1
      ^ state_4_4_49_lpi_3;
  assign state_4_8_sva_2_mx0w5 = xor_cse_673 ^ xor_cse_587 ^ xor_cse_702 ^ xor_cse_854;
  assign state_4_9_sva_2_mx0w5 = xor_cse_506 ^ xor_cse_469 ^ xor_cse_709 ^ state_4_4_9_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1 ^ state_1_1_63_32_lpi_4_23;
  assign xor_cse_859 = state_2_38_1_lpi_4 ^ state_0_38_lpi_6 ^ plaintext_63_32_sva_6
      ^ state_3_3_63_32_sva_6;
  assign xor_cse_858 = xor_cse_859 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_6 ^ Encrypt_Top_sbox_and_1_cse_38_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_38_sva_1;
  assign xor_cse_861 = plaintext_31_0_sva_10 ^ (state_4_3_31_0_sva_10 & plaintext_31_0_sva_10)
      ^ state_3_3_31_0_sva_10 ^ (plaintext_31_0_sva_10 & state_0_10_lpi_6);
  assign xor_cse_866 = state_2_38_1_lpi_4 ^ state_0_38_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_38_sva_1
      ^ xor_cse_588;
  assign xor_cse_867 = state_2_39_1_lpi_4 ^ state_0_39_lpi_6 ^ plaintext_63_32_sva_7
      ^ state_3_3_63_32_sva_7;
  assign xor_cse_868 = plaintext_31_0_sva_11 ^ (state_4_3_31_0_sva_11 & plaintext_31_0_sva_11)
      ^ state_3_3_31_0_sva_11 ^ (plaintext_31_0_sva_11 & state_0_11_lpi_6);
  assign xor_cse_871 = xor_cse_384 ^ Encrypt_Top_sbox_1_and_cse_30_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_30_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1;
  assign xor_cse_875 = state_1_1_63_32_lpi_4_13 ^ state_2_39_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_39_sva_1
      ^ state_3_39_lpi_3;
  assign xor_cse_878 = state_2_40_1_lpi_4 ^ state_0_40_lpi_6 ^ plaintext_63_32_sva_8
      ^ state_3_3_63_32_sva_8;
  assign xor_cse_877 = xor_cse_878 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_8 ^ Encrypt_Top_sbox_and_1_cse_40_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_40_sva_1;
  assign xor_cse_880 = plaintext_31_0_sva_12 ^ (state_4_3_31_0_sva_12 & plaintext_31_0_sva_12)
      ^ state_3_3_31_0_sva_12 ^ (plaintext_31_0_sva_12 & state_0_12_lpi_6);
  assign xor_cse_888 = state_2_41_1_lpi_4 ^ state_0_41_lpi_6 ^ plaintext_63_32_sva_9
      ^ state_3_3_63_32_sva_9;
  assign xor_cse_887 = xor_cse_888 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_9 ^ Encrypt_Top_sbox_and_1_cse_41_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_41_sva_1;
  assign xor_cse_890 = plaintext_31_0_sva_13 ^ (state_4_3_31_0_sva_13 & plaintext_31_0_sva_13)
      ^ state_3_3_31_0_sva_13 ^ (plaintext_31_0_sva_13 & state_0_13_lpi_6);
  assign xor_cse_895 = state_2_32_1_lpi_4 ^ state_0_32_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_32_sva_1
      ^ xor_cse_412;
  assign xor_cse_897 = state_1_1_63_32_lpi_4_15 ^ state_2_41_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_41_sva_1
      ^ state_3_41_lpi_3;
  assign xor_cse_899 = state_2_42_1_lpi_4 ^ state_0_42_lpi_6 ^ plaintext_63_32_sva_10
      ^ state_3_3_63_32_sva_10;
  assign xor_cse_900 = plaintext_31_0_sva_14 ^ (state_4_3_31_0_sva_14 & plaintext_31_0_sva_14)
      ^ state_3_3_31_0_sva_14 ^ (plaintext_31_0_sva_14 & state_0_14_lpi_6);
  assign xor_cse_905 = Encrypt_Top_sbox_2_and_2_cse_42_sva_1 ^ state_0_42_lpi_6;
  assign xor_cse_906 = state_2_33_1_lpi_4 ^ state_0_33_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_33_sva_1
      ^ xor_cse_425;
  assign xor_cse_910 = state_2_43_1_lpi_4 ^ state_0_43_lpi_6 ^ plaintext_63_32_sva_11
      ^ state_3_3_63_32_sva_11;
  assign xor_cse_909 = xor_cse_910 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_11 ^ Encrypt_Top_sbox_and_1_cse_43_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_43_sva_1;
  assign xor_cse_912 = plaintext_31_0_sva_15 ^ (state_4_3_31_0_sva_15 & plaintext_31_0_sva_15)
      ^ state_3_3_31_0_sva_15 ^ (plaintext_31_0_sva_15 & state_0_15_lpi_6);
  assign xor_cse_915 = state_2_43_1_lpi_4 ^ state_0_43_lpi_6 ^ xor_cse_151 ^ Encrypt_Top_sbox_1_and_1_cse_43_sva_1;
  assign xor_cse_920 = state_1_1_63_32_lpi_4_17 ^ state_2_43_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_43_sva_1
      ^ state_3_43_lpi_3;
  assign xor_cse_924 = state_2_44_1_lpi_4 ^ state_0_44_lpi_6 ^ plaintext_63_32_sva_12
      ^ state_3_3_63_32_sva_12;
  assign xor_cse_923 = xor_cse_924 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_12 ^ Encrypt_Top_sbox_and_1_cse_44_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_44_sva_1;
  assign xor_cse_926 = plaintext_31_0_sva_16 ^ (state_4_3_31_0_sva_16 & plaintext_31_0_sva_16)
      ^ state_3_3_31_0_sva_16 ^ (plaintext_31_0_sva_16 & state_0_16_lpi_6);
  assign xor_cse_927 = Encrypt_Top_sbox_and_1_cse_16_sva_1 ^ state_2_16_1_lpi_4 ^
      state_0_16_lpi_6;
  assign xor_cse_928 = state_0_44_lpi_6 ^ state_2_44_1_lpi_4 ^ Encrypt_Top_sbox_1_and_cse_16_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_16_sva_1;
  assign xor_cse_933 = plaintext_31_0_sva_17 ^ state_3_3_31_0_sva_17 ^ state_2_17_1_lpi_4
      ^ state_0_17_lpi_6;
  assign xor_cse_932 = xor_cse_933 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_17 ^ Encrypt_Top_sbox_and_1_cse_17_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_17_sva_1;
  assign xor_cse_935 = state_2_45_1_lpi_4 ^ state_0_45_lpi_6 ^ plaintext_63_32_sva_13
      ^ state_3_3_63_32_sva_13;
  assign xor_cse_936 = state_2_36_1_lpi_4 ^ state_0_36_lpi_6 ^ plaintext_63_32_sva_4
      ^ state_3_3_63_32_sva_4;
  assign xor_cse_943 = state_1_1_63_32_lpi_4_10 ^ state_2_36_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_36_sva_1
      ^ state_3_36_lpi_3;
  assign xor_cse_944 = state_1_1_63_32_lpi_4_19 ^ state_2_45_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_45_sva_1
      ^ state_3_45_lpi_3;
  assign xor_cse_948 = state_2_46_1_lpi_4 ^ state_0_46_lpi_6 ^ plaintext_63_32_sva_14
      ^ state_3_3_63_32_sva_14;
  assign xor_cse_947 = xor_cse_948 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_14 ^ Encrypt_Top_sbox_and_1_cse_46_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_46_sva_1;
  assign xor_cse_950 = state_2_37_1_lpi_4 ^ state_0_37_lpi_6 ^ plaintext_63_32_sva_5
      ^ state_3_3_63_32_sva_5;
  assign xor_cse_951 = plaintext_31_0_sva_18 ^ (state_4_3_31_0_sva_18 & plaintext_31_0_sva_18)
      ^ state_3_3_31_0_sva_18 ^ (plaintext_31_0_sva_18 & state_0_18_lpi_6);
  assign xor_cse_953 = Encrypt_Top_sbox_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_and_2_cse_37_sva_1;
  assign xor_cse_955 = state_2_46_1_lpi_4 ^ state_0_46_lpi_6 ^ state_0_37_lpi_6;
  assign xor_cse_958 = state_1_1_63_32_lpi_4_11 ^ state_2_37_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_37_sva_1
      ^ state_3_37_lpi_3;
  assign xor_cse_961 = state_2_47_1_lpi_4 ^ state_0_47_lpi_6 ^ plaintext_63_32_sva_15
      ^ state_3_3_63_32_sva_15;
  assign xor_cse_967 = state_1_1_63_32_lpi_4_20 ^ state_2_47_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_47_sva_1
      ^ state_3_47_lpi_3;
  assign xor_cse_970 = state_2_48_1_lpi_4 ^ state_0_48_lpi_6 ^ plaintext_63_32_sva_16
      ^ state_3_3_63_32_sva_16;
  assign xor_cse_977 = state_1_1_63_32_lpi_4_21 ^ state_2_48_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_48_sva_1
      ^ state_3_48_lpi_3;
  assign xor_cse_981 = state_2_49_1_lpi_4 ^ state_0_49_lpi_6 ^ plaintext_63_32_sva_17
      ^ state_3_3_63_32_sva_17;
  assign xor_cse_983 = xor_cse_290 ^ Encrypt_Top_sbox_1_and_1_cse_21_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_21_sva_1;
  assign xor_cse_985 = state_2_49_1_lpi_4 ^ state_0_49_lpi_6 ^ state_2_40_1_lpi_4
      ^ state_0_40_lpi_6;
  assign xor_cse_990 = state_2_50_1_lpi_4 ^ state_0_50_lpi_6 ^ plaintext_63_32_sva_18
      ^ state_3_3_63_32_sva_18;
  assign xor_cse_996 = state_1_1_63_32_lpi_4_23 ^ state_2_50_1_lpi_4 ^ Encrypt_Top_sbox_3_and_cse_50_sva_1
      ^ state_3_50_lpi_3;
  assign xor_cse_1000 = state_2_51_1_lpi_4 ^ state_0_51_lpi_6 ^ plaintext_63_32_sva_19
      ^ state_3_3_63_32_sva_19;
  assign xor_cse_1009 = state_2_52_1_lpi_4 ^ state_0_52_lpi_6 ^ plaintext_63_32_sva_20
      ^ state_3_3_63_32_sva_20;
  assign xor_cse_1016 = state_2_53_1_lpi_4 ^ state_0_53_lpi_6 ^ plaintext_63_32_sva_21
      ^ state_3_3_63_32_sva_21;
  assign xor_cse_1017 = Encrypt_Top_sbox_and_cse_63_32_sva_1_21 ^ Encrypt_Top_sbox_and_1_cse_53_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_53_sva_1;
  assign xor_cse_1018 = Encrypt_Top_sbox_1_and_1_cse_25_sva_1 ^ Encrypt_Top_sbox_1_and_cse_25_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1 ^ state_2_44_1_lpi_4;
  assign xor_cse_1021 = state_2_54_1_lpi_4 ^ state_0_54_lpi_6 ^ plaintext_63_32_sva_22
      ^ state_3_3_63_32_sva_22;
  assign xor_cse_1030 = state_2_55_1_lpi_4 ^ state_0_55_lpi_6 ^ plaintext_63_32_sva_23
      ^ state_3_3_63_32_sva_23;
  assign xor_cse_1031 = plaintext_31_0_sva_27 ^ (state_4_3_31_0_sva_27 & plaintext_31_0_sva_27)
      ^ state_3_3_31_0_sva_27 ^ (plaintext_31_0_sva_27 & state_0_27_lpi_6);
  assign xor_cse_1034 = xor_cse_343 ^ Encrypt_Top_sbox_1_and_cse_27_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_27_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_27_sva_1;
  assign xor_cse_1037 = state_2_55_1_lpi_4 ^ state_0_55_lpi_6;
  assign xor_cse_1041 = state_2_56_1_lpi_4 ^ state_0_56_lpi_6 ^ plaintext_63_32_sva_24
      ^ state_3_3_63_32_sva_24;
  assign xor_cse_1046 = state_2_56_1_lpi_4 ^ state_0_56_lpi_6;
  assign xor_cse_1050 = state_2_57_1_lpi_4 ^ state_0_57_lpi_6 ^ plaintext_63_32_sva_25
      ^ state_3_3_63_32_sva_25;
  assign xor_cse_1055 = state_2_57_1_lpi_4 ^ state_0_57_lpi_6;
  assign xor_cse_1059 = state_2_58_1_lpi_4 ^ state_0_58_lpi_6 ^ plaintext_63_32_sva_26
      ^ state_3_3_63_32_sva_26;
  assign xor_cse_1064 = state_2_58_1_lpi_4 ^ state_0_58_lpi_6;
  assign xor_cse_1068 = state_2_59_1_lpi_4 ^ state_0_59_lpi_6 ^ plaintext_63_32_sva_27
      ^ state_3_3_63_32_sva_27;
  assign xor_cse_1078 = plaintext_63_32_sva_28 ^ (state_4_3_63_32_sva_28 & plaintext_63_32_sva_28)
      ^ state_3_3_63_32_sva_28 ^ (plaintext_63_32_sva_28 & state_0_60_lpi_6);
  assign xor_cse_1077 = state_0_60_lpi_6 ^ state_2_60_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_60_sva_1
      ^ xor_cse_1078;
  assign xor_cse_1085 = state_2_60_1_lpi_4 ^ state_0_60_lpi_6;
  assign xor_cse_1087 = plaintext_63_32_sva_29 ^ (state_4_3_63_32_sva_29 & plaintext_63_32_sva_29)
      ^ state_3_3_63_32_sva_29 ^ (plaintext_63_32_sva_29 & state_0_61_lpi_6);
  assign xor_cse_1086 = state_0_61_lpi_6 ^ state_2_61_1_lpi_4 ^ Encrypt_Top_sbox_and_1_cse_61_sva_1
      ^ xor_cse_1087;
  assign xor_cse_1095 = state_2_61_1_lpi_4 ^ state_0_61_lpi_6;
  assign xor_cse_1097 = plaintext_63_32_sva_30 ^ (state_4_3_63_32_sva_30 & plaintext_63_32_sva_30)
      ^ state_3_3_63_32_sva_30 ^ (plaintext_63_32_sva_30 & state_0_62_lpi_6);
  assign xor_cse_1096 = state_2_62_1_lpi_4 ^ state_0_62_lpi_6 ^ Encrypt_Top_sbox_and_1_cse_62_sva_1
      ^ xor_cse_1097;
  assign xor_cse_1103 = state_2_63_1_lpi_4 ^ state_0_63_lpi_6 ^ plaintext_63_32_sva_31
      ^ state_3_3_63_32_sva_31;
  assign xor_cse_1108 = state_2_63_1_lpi_4 ^ state_0_63_lpi_6;
  assign state_0_8_sva_3_mx0w5 = xor_cse_1034 ^ xor_cse_159 ^ xor_cse_59 ^ Encrypt_Top_sbox_1_and_1_cse_8_sva_1
      ^ state_2_8_1_lpi_4 ^ state_0_8_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_36_sva_1
      ^ state_2_36_1_lpi_4 ^ state_0_36_lpi_6;
  assign state_0_9_sva_3_mx0w5 = xor_cse_356 ^ xor_cse_170 ^ xor_cse_74 ^ Encrypt_Top_sbox_1_and_1_cse_9_sva_1
      ^ state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1
      ^ state_2_37_1_lpi_4 ^ state_0_37_lpi_6;
  assign xor_cse_1134 = xor_cse_102 ^ state_0_3_lpi_6 ^ state_2_58_1_lpi_4 ^ state_0_58_lpi_6
      ^ state_0_39_lpi_6 ^ state_2_3_1_lpi_4;
  assign xor_cse_1144 = state_2_4_1_lpi_4 ^ state_0_4_lpi_6 ^ state_2_40_1_lpi_4
      ^ state_0_40_lpi_6;
  assign xor_cse_1162 = state_2_8_1_lpi_4 ^ state_0_8_lpi_6 ^ state_3_3_31_0_sva_8
      ^ plaintext_31_0_sva_8;
  assign xor_cse_1161 = xor_cse_1162 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_8 ^ Encrypt_Top_sbox_and_1_cse_8_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_8_sva_1;
  assign xor_cse_1167 = state_2_8_1_lpi_4 ^ state_0_8_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_8_sva_1
      ^ xor_cse_587;
  assign xor_cse_1172 = state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ state_3_3_31_0_sva_9
      ^ plaintext_31_0_sva_9;
  assign xor_cse_1171 = xor_cse_1172 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_9 ^ Encrypt_Top_sbox_and_1_cse_9_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_9_sva_1;
  assign xor_cse_1187 = state_2_12_1_lpi_4 ^ state_0_12_lpi_6;
  assign xor_cse_1188 = xor_cse_102 ^ state_0_3_lpi_6 ^ state_2_3_1_lpi_4 ^ xor_cse_204;
  assign xor_cse_1193 = state_2_13_1_lpi_4 ^ state_0_13_lpi_6;
  assign xor_cse_1293 = state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6])
      ^ (state_4_3_31_0_sva_6 & state_3_3_31_0_sva_6) ^ state_4_3_31_0_sva_6;
  assign xor_cse_1299 = state_4_4_17_lpi_3 ^ Encrypt_Top_sbox_2_and_656 ^ Encrypt_Top_sbox_2_and_658
      ^ Encrypt_Top_sbox_2_and_600;
  assign xor_cse_1300 = xor_cse_178 ^ Encrypt_Top_sbox_2_and_602 ^ state_4_4_10_lpi_3
      ^ xor_cse_196;
  assign state_3_0_sva_3_mx0w6 = xor_cse_252 ^ xor_cse_197 ^ xor_cse_1299 ^ xor_cse_1300;
  assign xor_cse_1301 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]) ^ Encrypt_Top_sbox_1_and_768
      ^ state_4_4_6_lpi_3 ^ state_1_1_31_0_lpi_4_6;
  assign state_2_0_1_sva_4 = ~(xor_cse_806 ^ xor_cse_813 ^ xor_cse_1301 ^ state_2_0_1_lpi_4
      ^ state_2_1_1_lpi_4 ^ state_2_6_1_lpi_4);
  assign xor_cse_1303 = state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7])
      ^ (state_4_3_31_0_sva_7 & state_3_3_31_0_sva_7) ^ state_4_3_31_0_sva_7;
  assign xor_cse_1306 = state_2_7_1_lpi_4 ^ Encrypt_Top_sbox_1_and_770 ^ state_4_4_7_lpi_3
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7]);
  assign xor_cse_1309 = state_4_4_18_lpi_3 ^ Encrypt_Top_sbox_2_and_664 ^ Encrypt_Top_sbox_2_and_666
      ^ Encrypt_Top_sbox_2_and_608;
  assign xor_cse_1310 = Encrypt_Top_sbox_2_and_610 ^ state_4_4_11_lpi_3;
  assign state_3_1_sva_3_mx0w6 = xor_cse_206 ^ xor_cse_189 ^ xor_cse_263 ^ xor_cse_207
      ^ xor_cse_1309 ^ xor_cse_1310;
  assign xor_cse_1311 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]) ^ Encrypt_Top_sbox_1_and_770
      ^ state_4_4_7_lpi_3 ^ state_1_1_31_0_lpi_4_7;
  assign state_2_1_1_sva_4 = ~(xor_cse_813 ^ xor_cse_821 ^ xor_cse_1311 ^ state_2_1_1_lpi_4
      ^ state_2_2_1_lpi_4 ^ state_2_7_1_lpi_4);
  assign xor_cse_1317 = xor_cse_343 ^ (state_4_4_27_lpi_3 & state_0_27_lpi_6) ^ (state_3_27_lpi_3
      & state_0_27_lpi_6) ^ state_4_4_27_lpi_3;
  assign state_3_10_sva_2_mx0w6 = xor_cse_1317 ^ xor_cse_178 ^ xor_cse_282 ^ Encrypt_Top_sbox_2_and_600
      ^ Encrypt_Top_sbox_2_and_602 ^ state_4_4_10_lpi_3 ^ Encrypt_Top_sbox_2_and_680
      ^ Encrypt_Top_sbox_2_and_682 ^ state_4_4_20_lpi_3;
  assign state_2_2_1_sva_4 = ~(xor_cse_821 ^ xor_cse_826 ^ xor_cse_850 ^ state_2_2_1_lpi_4
      ^ state_2_3_1_lpi_4);
  assign xor_cse_1324 = state_4_4_28_lpi_3 ^ (state_4_4_28_lpi_3 & state_0_28_lpi_6)
      ^ (state_3_28_lpi_3 & state_0_28_lpi_6) ^ xor_cse_357;
  assign xor_cse_1325 = xor_cse_290 ^ Encrypt_Top_sbox_2_and_688 ^ Encrypt_Top_sbox_2_and_690
      ^ state_4_4_21_lpi_3;
  assign state_3_11_sva_2_mx0w6 = xor_cse_1324 ^ xor_cse_1325 ^ xor_cse_189 ^ Encrypt_Top_sbox_2_and_608
      ^ Encrypt_Top_sbox_2_and_610 ^ state_4_4_11_lpi_3;
  assign state_2_3_1_sva_4 = ~(xor_cse_826 ^ xor_cse_833 ^ xor_cse_851 ^ state_2_3_1_lpi_4
      ^ state_2_4_1_lpi_4);
  assign xor_cse_1332 = xor_cse_299 ^ Encrypt_Top_sbox_2_and_698 ^ state_4_4_22_lpi_3
      ^ Encrypt_Top_sbox_2_and_696;
  assign state_3_12_sva_2_mx0w6 = xor_cse_1332 ^ xor_cse_204 ^ xor_cse_369 ^ Encrypt_Top_sbox_2_and_616
      ^ Encrypt_Top_sbox_2_and_618 ^ state_4_4_12_lpi_3 ^ Encrypt_Top_sbox_2_and_752
      ^ Encrypt_Top_sbox_2_and_754 ^ state_4_4_29_lpi_3;
  assign state_2_4_1_sva_4 = ~(xor_cse_465 ^ xor_cse_833 ^ xor_cse_839 ^ state_2_4_1_lpi_4
      ^ state_2_5_1_lpi_4);
  assign xor_cse_1341 = xor_cse_384 ^ (state_4_4_30_lpi_3 & state_0_30_lpi_6) ^ (state_3_30_lpi_3
      & state_0_30_lpi_6) ^ state_4_4_30_lpi_3;
  assign state_3_13_sva_2_mx0w6 = xor_cse_1341 ^ xor_cse_211 ^ xor_cse_308 ^ Encrypt_Top_sbox_2_and_624
      ^ Encrypt_Top_sbox_2_and_704 ^ Encrypt_Top_sbox_2_and_706 ^ Encrypt_Top_sbox_2_and_626
      ^ state_4_4_13_lpi_3 ^ state_4_4_23_lpi_3;
  assign state_2_5_1_sva_4 = ~(xor_cse_839 ^ xor_cse_1301 ^ xor_cse_466 ^ state_2_5_1_lpi_4
      ^ state_2_6_1_lpi_4);
  assign xor_cse_1350 = xor_cse_316 ^ (state_4_4_24_lpi_3 & state_0_24_lpi_6) ^ (state_3_24_lpi_3
      & state_0_24_lpi_6) ^ state_4_4_24_lpi_3;
  assign xor_cse_1351 = xor_cse_394 ^ (state_4_4_31_lpi_3 & state_0_31_lpi_6) ^ (state_3_31_lpi_3
      & state_0_31_lpi_6) ^ state_4_4_31_lpi_3;
  assign state_3_14_sva_2_mx0w6 = xor_cse_1350 ^ xor_cse_1351 ^ xor_cse_221 ^ Encrypt_Top_sbox_2_and_632
      ^ Encrypt_Top_sbox_2_and_634 ^ state_4_4_14_lpi_3;
  assign state_2_6_1_sva_4 = ~(xor_cse_1301 ^ xor_cse_1311 ^ xor_cse_477 ^ state_2_6_1_lpi_4
      ^ state_2_7_1_lpi_4);
  assign xor_cse_1357 = xor_cse_325 ^ (state_4_4_25_lpi_3 & state_0_25_lpi_6) ^ (state_3_25_lpi_3
      & state_0_25_lpi_6) ^ state_4_4_25_lpi_3;
  assign xor_cse_1358 = state_1_1_31_0_lpi_4_8 ^ xor_cse_11 ^ Encrypt_Top_sbox_2_and_764
      ^ Encrypt_Top_sbox_2_and_766;
  assign xor_cse_1360 = Encrypt_Top_sbox_2_and_640 ^ Encrypt_Top_sbox_2_and_642 ^
      state_4_4_15_lpi_3;
  assign state_3_15_sva_3_mx0w6 = xor_cse_1357 ^ xor_cse_1358 ^ xor_cse_231 ^ xor_cse_1360;
  assign state_2_7_1_sva_4 = ~(state_2_7_1_lpi_4 ^ xor_cse_1311 ^ xor_cse_850 ^ xor_cse_488);
  assign xor_cse_1361 = xor_cse_430 ^ Encrypt_Top_sbox_and_1_cse_6_sva_1 ^ plaintext_31_0_sva_6
      ^ state_4_3_31_0_sva_6;
  assign xor_cse_1363 = INIT_P12_INIT_P12_xor_2_psp_sva_1 & state_3_3_31_0_sva_6;
  assign xor_cse_1364 = state_3_3_31_0_sva_6 & plaintext_31_0_sva_6;
  assign xor_cse_1366 = plaintext_31_0_sva_28 ^ state_3_3_31_0_sva_28 ^ state_4_3_31_0_sva_28
      ^ state_2_28_1_lpi_4;
  assign xor_cse_1367 = plaintext_31_0_sva_31 ^ state_3_3_31_0_sva_31 ^ state_4_3_31_0_sva_31
      ^ state_2_31_1_lpi_4;
  assign xor_cse_1368 = (state_2_31_1_lpi_4 & state_3_3_31_0_sva_31) ^ (state_3_3_31_0_sva_31
      & plaintext_31_0_sva_31) ^ Encrypt_Top_sbox_and_1_cse_31_sva_1 ^ state_0_31_lpi_6;
  assign xor_cse_1371 = (state_2_28_1_lpi_4 & state_3_3_31_0_sva_28) ^ (state_3_3_31_0_sva_28
      & plaintext_31_0_sva_28) ^ Encrypt_Top_sbox_and_1_cse_28_sva_1 ^ state_0_28_lpi_6;
  assign state_1_1_31_0_sva_1_31_1 = xor_cse_1361 ^ xor_cse_1363 ^ xor_cse_1364 ^
      xor_cse_1366 ^ xor_cse_1367 ^ xor_cse_1368 ^ xor_cse_1371;
  assign xor_cse_1375 = plaintext_63_32_sva_29 ^ state_3_3_63_32_sva_29 ^ state_4_3_63_32_sva_29
      ^ state_2_61_1_lpi_4;
  assign xor_cse_1374 = state_0_61_lpi_6 ^ xor_cse_1375 ^ (state_2_61_1_lpi_4 & state_3_3_63_32_sva_29)
      ^ (state_3_3_63_32_sva_29 & plaintext_63_32_sva_29);
  assign xor_cse_1378 = xor_cse_352 ^ Encrypt_Top_sbox_and_1_cse_0_sva_1 ^ plaintext_31_0_sva_0
      ^ state_4_3_31_0_sva_0;
  assign xor_cse_1381 = INIT_P12_INIT_P12_xor_8_psp_sva_1 & state_3_3_31_0_sva_0;
  assign xor_cse_1382 = state_3_3_31_0_sva_0 & plaintext_31_0_sva_0;
  assign xor_cse_1384 = state_2_39_1_lpi_4 & state_3_3_63_32_sva_7;
  assign xor_cse_1385 = state_3_3_63_32_sva_7 & plaintext_63_32_sva_7;
  assign state_1_1_31_0_sva_1_0_1 = xor_cse_1374 ^ xor_cse_1378 ^ xor_cse_867 ^ xor_cse_1381
      ^ xor_cse_1382 ^ Encrypt_Top_sbox_and_1_cse_61_sva_1 ^ state_4_3_63_32_sva_7
      ^ xor_cse_1384 ^ xor_cse_1385 ^ Encrypt_Top_sbox_and_1_cse_39_sva_1;
  assign xor_cse_1386 = xor_cse_417 ^ Encrypt_Top_sbox_and_1_cse_5_sva_1 ^ plaintext_31_0_sva_5
      ^ state_4_3_31_0_sva_5;
  assign xor_cse_1388 = INIT_P12_INIT_P12_xor_3_psp_sva_1 & state_3_3_31_0_sva_5;
  assign xor_cse_1389 = state_3_3_31_0_sva_5 & plaintext_31_0_sva_5;
  assign xor_cse_1391 = plaintext_31_0_sva_30 ^ state_3_3_31_0_sva_30 ^ state_4_3_31_0_sva_30
      ^ state_2_30_1_lpi_4;
  assign xor_cse_1392 = plaintext_31_0_sva_27 ^ state_3_3_31_0_sva_27 ^ state_4_3_31_0_sva_27
      ^ state_2_27_1_lpi_4;
  assign xor_cse_1393 = (state_2_30_1_lpi_4 & state_3_3_31_0_sva_30) ^ (state_3_3_31_0_sva_30
      & plaintext_31_0_sva_30) ^ Encrypt_Top_sbox_and_1_cse_30_sva_1 ^ state_0_30_lpi_6;
  assign xor_cse_1396 = (state_2_27_1_lpi_4 & state_3_3_31_0_sva_27) ^ (state_3_3_31_0_sva_27
      & plaintext_31_0_sva_27) ^ Encrypt_Top_sbox_and_1_cse_27_sva_1 ^ state_0_27_lpi_6;
  assign state_1_1_31_0_sva_1_30_1 = xor_cse_1386 ^ xor_cse_1388 ^ xor_cse_1389 ^
      xor_cse_1391 ^ xor_cse_1392 ^ xor_cse_1393 ^ xor_cse_1396;
  assign xor_cse_1400 = plaintext_63_32_sva_30 ^ state_3_3_63_32_sva_30 ^ state_4_3_63_32_sva_30
      ^ state_2_62_1_lpi_4;
  assign xor_cse_1399 = state_0_62_lpi_6 ^ xor_cse_1400 ^ (state_2_62_1_lpi_4 & state_3_3_63_32_sva_30)
      ^ (state_3_3_63_32_sva_30 & plaintext_63_32_sva_30);
  assign xor_cse_1403 = xor_cse_878 ^ state_4_3_63_32_sva_8 ^ (state_2_40_1_lpi_4
      & state_3_3_63_32_sva_8) ^ (state_3_3_63_32_sva_8 & plaintext_63_32_sva_8);
  assign xor_cse_1406 = xor_cse_364 ^ Encrypt_Top_sbox_and_1_cse_1_sva_1 ^ plaintext_31_0_sva_1
      ^ state_4_3_31_0_sva_1;
  assign xor_cse_1408 = INIT_P12_INIT_P12_xor_7_psp_sva_1 & state_3_3_31_0_sva_1;
  assign xor_cse_1409 = state_3_3_31_0_sva_1 & plaintext_31_0_sva_1;
  assign state_1_1_31_0_sva_1_1_1 = xor_cse_1399 ^ xor_cse_1403 ^ xor_cse_1406 ^
      xor_cse_1408 ^ xor_cse_1409 ^ Encrypt_Top_sbox_and_1_cse_62_sva_1 ^ Encrypt_Top_sbox_and_1_cse_40_sva_1;
  assign xor_cse_1410 = xor_cse_405 ^ Encrypt_Top_sbox_and_1_cse_4_sva_1 ^ plaintext_31_0_sva_4
      ^ state_4_3_31_0_sva_4;
  assign xor_cse_1412 = INIT_P12_INIT_P12_xor_4_psp_sva_1 & state_3_3_31_0_sva_4;
  assign xor_cse_1413 = state_3_3_31_0_sva_4 & plaintext_31_0_sva_4;
  assign xor_cse_1415 = plaintext_31_0_sva_29 ^ state_3_3_31_0_sva_29 ^ state_4_3_31_0_sva_29
      ^ state_2_29_1_lpi_4;
  assign xor_cse_1416 = plaintext_31_0_sva_26 ^ state_3_3_31_0_sva_26 ^ state_4_3_31_0_sva_26
      ^ state_2_26_1_lpi_4;
  assign xor_cse_1418 = state_2_29_1_lpi_4 & state_3_3_31_0_sva_29;
  assign xor_cse_1419 = state_3_3_31_0_sva_29 & plaintext_31_0_sva_29;
  assign xor_cse_1417 = xor_cse_1418 ^ xor_cse_1419 ^ Encrypt_Top_sbox_and_1_cse_29_sva_1
      ^ state_0_29_lpi_6;
  assign xor_cse_1420 = (state_2_26_1_lpi_4 & state_3_3_31_0_sva_26) ^ (state_3_3_31_0_sva_26
      & plaintext_31_0_sva_26) ^ Encrypt_Top_sbox_and_1_cse_26_sva_1 ^ state_0_26_lpi_6;
  assign state_1_1_31_0_sva_1_29_1 = xor_cse_1410 ^ xor_cse_1412 ^ xor_cse_1413 ^
      xor_cse_1415 ^ xor_cse_1416 ^ xor_cse_1417 ^ xor_cse_1420;
  assign xor_cse_1423 = xor_cse_888 ^ state_4_3_63_32_sva_9 ^ (state_2_41_1_lpi_4
      & state_3_3_63_32_sva_9) ^ (state_3_3_63_32_sva_9 & plaintext_63_32_sva_9);
  assign xor_cse_1426 = xor_cse_377 ^ Encrypt_Top_sbox_and_1_cse_2_sva_1 ^ plaintext_31_0_sva_2
      ^ state_4_3_31_0_sva_2;
  assign xor_cse_1429 = INIT_P12_INIT_P12_xor_6_psp_sva_1 & state_3_3_31_0_sva_2;
  assign xor_cse_1430 = state_3_3_31_0_sva_2 & plaintext_31_0_sva_2;
  assign xor_cse_1431 = state_2_63_1_lpi_4 & state_3_3_63_32_sva_31;
  assign xor_cse_1433 = state_3_3_63_32_sva_31 & plaintext_63_32_sva_31;
  assign state_1_1_31_0_sva_1_2_1 = xor_cse_1423 ^ xor_cse_1426 ^ xor_cse_1103 ^
      xor_cse_1429 ^ xor_cse_1430 ^ state_4_3_63_32_sva_31 ^ xor_cse_1431 ^ xor_cse_1433
      ^ Encrypt_Top_sbox_and_1_cse_63_sva_1 ^ Encrypt_Top_sbox_and_1_cse_41_sva_1;
  assign xor_cse_1434 = xor_cse_389 ^ Encrypt_Top_sbox_and_1_cse_3_sva_1 ^ plaintext_31_0_sva_3
      ^ state_4_3_31_0_sva_3;
  assign xor_cse_1436 = INIT_P12_INIT_P12_xor_5_psp_sva_1 & state_3_3_31_0_sva_3;
  assign xor_cse_1437 = state_3_3_31_0_sva_3 & plaintext_31_0_sva_3;
  assign xor_cse_1439 = plaintext_31_0_sva_25 ^ state_3_3_31_0_sva_25 ^ state_4_3_31_0_sva_25
      ^ state_2_25_1_lpi_4;
  assign xor_cse_1441 = (state_2_25_1_lpi_4 & state_3_3_31_0_sva_25) ^ (state_3_3_31_0_sva_25
      & plaintext_31_0_sva_25) ^ Encrypt_Top_sbox_and_1_cse_25_sva_1 ^ state_0_25_lpi_6;
  assign state_1_1_31_0_sva_1_28_1 = xor_cse_1434 ^ xor_cse_1436 ^ xor_cse_1437 ^
      xor_cse_1366 ^ xor_cse_1439 ^ xor_cse_1371 ^ xor_cse_1441;
  assign xor_cse_1446 = state_4_3_63_32_sva_10 ^ (state_2_42_1_lpi_4 & state_3_3_63_32_sva_10)
      ^ (state_3_3_63_32_sva_10 & plaintext_63_32_sva_10) ^ Encrypt_Top_sbox_and_1_cse_42_sva_1;
  assign state_1_1_31_0_sva_1_3_1 = xor_cse_1378 ^ xor_cse_1434 ^ xor_cse_899 ^ xor_cse_1436
      ^ xor_cse_1437 ^ xor_cse_1381 ^ xor_cse_1382 ^ xor_cse_1446;
  assign xor_cse_1451 = plaintext_31_0_sva_24 ^ state_3_3_31_0_sva_24 ^ state_4_3_31_0_sva_24
      ^ state_2_24_1_lpi_4;
  assign xor_cse_1454 = state_2_24_1_lpi_4 & state_3_3_31_0_sva_24;
  assign xor_cse_1455 = state_3_3_31_0_sva_24 & plaintext_31_0_sva_24;
  assign xor_cse_1453 = xor_cse_1454 ^ xor_cse_1455 ^ Encrypt_Top_sbox_and_1_cse_24_sva_1
      ^ state_0_24_lpi_6;
  assign state_1_1_31_0_sva_1_27_1 = xor_cse_1426 ^ xor_cse_1429 ^ xor_cse_1430 ^
      xor_cse_1451 ^ xor_cse_1392 ^ xor_cse_1396 ^ xor_cse_1453;
  assign xor_cse_1456 = xor_cse_910 ^ state_4_3_63_32_sva_11 ^ (state_2_43_1_lpi_4
      & state_3_3_63_32_sva_11) ^ (state_3_3_63_32_sva_11 & plaintext_63_32_sva_11);
  assign state_1_1_31_0_sva_1_4_1 = xor_cse_1456 ^ xor_cse_1406 ^ xor_cse_1410 ^
      Encrypt_Top_sbox_and_1_cse_43_sva_1 ^ xor_cse_1412 ^ xor_cse_1413 ^ xor_cse_1408
      ^ xor_cse_1409;
  assign xor_cse_1463 = plaintext_31_0_sva_23 ^ state_3_3_31_0_sva_23 ^ state_4_3_31_0_sva_23
      ^ state_2_23_1_lpi_4;
  assign xor_cse_1465 = (state_2_23_1_lpi_4 & state_3_3_31_0_sva_23) ^ (state_3_3_31_0_sva_23
      & plaintext_31_0_sva_23) ^ Encrypt_Top_sbox_and_1_cse_23_sva_1 ^ state_0_23_lpi_6;
  assign state_1_1_31_0_sva_1_26_1 = xor_cse_1406 ^ xor_cse_1408 ^ xor_cse_1409 ^
      xor_cse_1463 ^ xor_cse_1416 ^ xor_cse_1420 ^ xor_cse_1465;
  assign xor_cse_1468 = xor_cse_924 ^ state_4_3_63_32_sva_12 ^ (state_2_44_1_lpi_4
      & state_3_3_63_32_sva_12) ^ (state_3_3_63_32_sva_12 & plaintext_63_32_sva_12);
  assign state_1_1_31_0_sva_1_5_1 = xor_cse_1468 ^ xor_cse_1426 ^ xor_cse_1386 ^
      Encrypt_Top_sbox_and_1_cse_44_sva_1 ^ xor_cse_1388 ^ xor_cse_1389 ^ xor_cse_1429
      ^ xor_cse_1430;
  assign xor_cse_1475 = plaintext_31_0_sva_22 ^ state_3_3_31_0_sva_22 ^ state_4_3_31_0_sva_22
      ^ state_2_22_1_lpi_4;
  assign xor_cse_1478 = state_2_22_1_lpi_4 & state_3_3_31_0_sva_22;
  assign xor_cse_1479 = state_3_3_31_0_sva_22 & plaintext_31_0_sva_22;
  assign xor_cse_1477 = xor_cse_1478 ^ xor_cse_1479 ^ Encrypt_Top_sbox_and_1_cse_22_sva_1
      ^ state_0_22_lpi_6;
  assign state_1_1_31_0_sva_1_25_1 = xor_cse_1378 ^ xor_cse_1381 ^ xor_cse_1382 ^
      xor_cse_1475 ^ xor_cse_1439 ^ xor_cse_1441 ^ xor_cse_1477;
  assign xor_cse_1482 = state_4_3_63_32_sva_13 ^ (state_2_45_1_lpi_4 & state_3_3_63_32_sva_13)
      ^ (state_3_3_63_32_sva_13 & plaintext_63_32_sva_13) ^ Encrypt_Top_sbox_and_1_cse_45_sva_1;
  assign state_1_1_31_0_sva_1_6_1 = xor_cse_1434 ^ xor_cse_1361 ^ xor_cse_935 ^ xor_cse_1363
      ^ xor_cse_1364 ^ xor_cse_1436 ^ xor_cse_1437 ^ xor_cse_1482;
  assign xor_cse_1485 = plaintext_31_0_sva_21 ^ state_3_3_31_0_sva_21 ^ state_4_3_31_0_sva_21
      ^ state_2_21_1_lpi_4;
  assign xor_cse_1488 = state_2_21_1_lpi_4 & state_3_3_31_0_sva_21;
  assign xor_cse_1489 = state_3_3_31_0_sva_21 & plaintext_31_0_sva_21;
  assign xor_cse_1487 = xor_cse_1488 ^ xor_cse_1489 ^ Encrypt_Top_sbox_and_1_cse_21_sva_1
      ^ state_0_21_lpi_6;
  assign xor_cse_1490 = state_4_3_63_32_sva_31 ^ xor_cse_1431 ^ xor_cse_1433 ^ Encrypt_Top_sbox_and_1_cse_63_sva_1;
  assign state_1_1_31_0_sva_1_24_1 = xor_cse_1103 ^ xor_cse_1485 ^ xor_cse_1451 ^
      xor_cse_1453 ^ xor_cse_1487 ^ xor_cse_1490;
  assign xor_cse_1491 = xor_cse_444 ^ Encrypt_Top_sbox_and_1_cse_7_sva_1 ^ plaintext_31_0_sva_7
      ^ state_4_3_31_0_sva_7;
  assign xor_cse_1492 = xor_cse_948 ^ state_4_3_63_32_sva_14 ^ (state_2_46_1_lpi_4
      & state_3_3_63_32_sva_14) ^ (state_3_3_63_32_sva_14 & plaintext_63_32_sva_14);
  assign xor_cse_1497 = INIT_P12_INIT_P12_xor_1_psp_sva_1 & state_3_3_31_0_sva_7;
  assign xor_cse_1498 = state_3_3_31_0_sva_7 & plaintext_31_0_sva_7;
  assign state_1_1_31_0_sva_1_7_1 = xor_cse_1491 ^ xor_cse_1492 ^ xor_cse_1410 ^
      Encrypt_Top_sbox_and_1_cse_46_sva_1 ^ xor_cse_1497 ^ xor_cse_1498 ^ xor_cse_1412
      ^ xor_cse_1413;
  assign xor_cse_1499 = (state_2_20_1_lpi_4 & state_3_3_31_0_sva_20) ^ (state_3_3_31_0_sva_20
      & plaintext_31_0_sva_20) ^ Encrypt_Top_sbox_and_1_cse_20_sva_1 ^ state_0_20_lpi_6;
  assign xor_cse_1503 = plaintext_31_0_sva_20 ^ state_3_3_31_0_sva_20 ^ state_4_3_31_0_sva_20
      ^ state_2_20_1_lpi_4;
  assign state_1_1_31_0_sva_1_23_1 = xor_cse_1399 ^ xor_cse_1499 ^ Encrypt_Top_sbox_and_1_cse_62_sva_1
      ^ xor_cse_1503 ^ xor_cse_1463 ^ xor_cse_1465;
  assign xor_cse_1505 = xor_cse_1162 ^ state_4_3_31_0_sva_8 ^ (state_2_8_1_lpi_4
      & state_3_3_31_0_sva_8) ^ (state_3_3_31_0_sva_8 & plaintext_31_0_sva_8);
  assign xor_cse_1511 = state_2_47_1_lpi_4 & state_3_3_63_32_sva_15;
  assign xor_cse_1512 = state_3_3_63_32_sva_15 & plaintext_63_32_sva_15;
  assign state_1_1_31_0_sva_1_8_1 = xor_cse_1505 ^ xor_cse_1386 ^ xor_cse_961 ^ Encrypt_Top_sbox_and_1_cse_8_sva_1
      ^ xor_cse_1388 ^ xor_cse_1389 ^ state_4_3_63_32_sva_15 ^ xor_cse_1511 ^ xor_cse_1512
      ^ Encrypt_Top_sbox_and_1_cse_47_sva_1;
  assign xor_cse_1514 = state_2_19_1_lpi_4 & state_3_3_31_0_sva_19;
  assign xor_cse_1515 = state_3_3_31_0_sva_19 & plaintext_31_0_sva_19;
  assign xor_cse_1513 = xor_cse_1514 ^ xor_cse_1515 ^ Encrypt_Top_sbox_and_1_cse_19_sva_1
      ^ state_0_19_lpi_6;
  assign xor_cse_1517 = plaintext_31_0_sva_19 ^ state_3_3_31_0_sva_19 ^ state_4_3_31_0_sva_19
      ^ state_2_19_1_lpi_4;
  assign state_1_1_31_0_sva_1_22_1 = xor_cse_1374 ^ xor_cse_1513 ^ Encrypt_Top_sbox_and_1_cse_61_sva_1
      ^ xor_cse_1517 ^ xor_cse_1475 ^ xor_cse_1477;
  assign xor_cse_1519 = xor_cse_1172 ^ state_4_3_31_0_sva_9 ^ (state_2_9_1_lpi_4
      & state_3_3_31_0_sva_9) ^ (state_3_3_31_0_sva_9 & plaintext_31_0_sva_9);
  assign xor_cse_1525 = state_2_48_1_lpi_4 & state_3_3_63_32_sva_16;
  assign xor_cse_1526 = state_3_3_63_32_sva_16 & plaintext_63_32_sva_16;
  assign state_1_1_31_0_sva_1_9_1 = xor_cse_1519 ^ xor_cse_1361 ^ xor_cse_970 ^ Encrypt_Top_sbox_and_1_cse_9_sva_1
      ^ xor_cse_1363 ^ xor_cse_1364 ^ state_4_3_63_32_sva_16 ^ xor_cse_1525 ^ xor_cse_1526
      ^ Encrypt_Top_sbox_and_1_cse_48_sva_1;
  assign xor_cse_1528 = plaintext_63_32_sva_28 ^ state_3_3_63_32_sva_28 ^ state_4_3_63_32_sva_28
      ^ state_2_60_1_lpi_4;
  assign xor_cse_1527 = state_0_60_lpi_6 ^ xor_cse_1528 ^ (state_2_60_1_lpi_4 & state_3_3_63_32_sva_28)
      ^ (state_3_3_63_32_sva_28 & plaintext_63_32_sva_28);
  assign xor_cse_1532 = state_2_18_1_lpi_4 & state_3_3_31_0_sva_18;
  assign xor_cse_1533 = state_3_3_31_0_sva_18 & plaintext_31_0_sva_18;
  assign xor_cse_1531 = xor_cse_1532 ^ xor_cse_1533 ^ Encrypt_Top_sbox_and_1_cse_18_sva_1
      ^ state_0_18_lpi_6;
  assign xor_cse_1535 = plaintext_31_0_sva_18 ^ state_3_3_31_0_sva_18 ^ state_4_3_31_0_sva_18
      ^ state_2_18_1_lpi_4;
  assign state_1_1_31_0_sva_1_21_1 = xor_cse_1527 ^ xor_cse_1531 ^ Encrypt_Top_sbox_and_1_cse_60_sva_1
      ^ xor_cse_1485 ^ xor_cse_1535 ^ xor_cse_1487;
  assign xor_cse_1538 = state_3_3_63_32_sva_17 & plaintext_63_32_sva_17;
  assign xor_cse_1540 = plaintext_31_0_sva_10 ^ state_3_3_31_0_sva_10 ^ state_4_3_31_0_sva_10
      ^ state_2_10_1_lpi_4;
  assign xor_cse_1542 = state_2_10_1_lpi_4 & state_3_3_31_0_sva_10;
  assign xor_cse_1543 = state_3_3_31_0_sva_10 & plaintext_31_0_sva_10;
  assign xor_cse_1541 = xor_cse_1542 ^ xor_cse_1543 ^ Encrypt_Top_sbox_and_1_cse_10_sva_1
      ^ state_0_10_lpi_6;
  assign xor_cse_1545 = state_2_49_1_lpi_4 & state_3_3_63_32_sva_17;
  assign state_1_1_31_0_sva_1_10_1 = xor_cse_1491 ^ xor_cse_1538 ^ Encrypt_Top_sbox_and_1_cse_49_sva_1
      ^ xor_cse_981 ^ xor_cse_1540 ^ xor_cse_1541 ^ xor_cse_1497 ^ xor_cse_1498 ^
      state_4_3_63_32_sva_17 ^ xor_cse_1545;
  assign xor_cse_1546 = xor_cse_933 ^ state_4_3_31_0_sva_17 ^ (state_2_17_1_lpi_4
      & state_3_3_31_0_sva_17) ^ (state_3_3_31_0_sva_17 & plaintext_31_0_sva_17);
  assign xor_cse_1550 = state_2_59_1_lpi_4 & state_3_3_63_32_sva_27;
  assign xor_cse_1551 = state_3_3_63_32_sva_27 & plaintext_63_32_sva_27;
  assign state_1_1_31_0_sva_1_20_1 = xor_cse_1546 ^ Encrypt_Top_sbox_and_1_cse_17_sva_1
      ^ state_4_3_63_32_sva_27 ^ xor_cse_1550 ^ xor_cse_1551 ^ Encrypt_Top_sbox_and_1_cse_59_sva_1
      ^ xor_cse_1068 ^ xor_cse_1503 ^ xor_cse_1499;
  assign xor_cse_1555 = state_2_50_1_lpi_4 & state_3_3_63_32_sva_18;
  assign xor_cse_1556 = state_3_3_63_32_sva_18 & plaintext_63_32_sva_18;
  assign xor_cse_1558 = plaintext_31_0_sva_11 ^ state_3_3_31_0_sva_11 ^ state_4_3_31_0_sva_11
      ^ state_2_11_1_lpi_4;
  assign xor_cse_1559 = (state_2_11_1_lpi_4 & state_3_3_31_0_sva_11) ^ (state_3_3_31_0_sva_11
      & plaintext_31_0_sva_11) ^ Encrypt_Top_sbox_and_1_cse_11_sva_1 ^ state_0_11_lpi_6;
  assign state_1_1_31_0_sva_1_11_1 = xor_cse_1505 ^ Encrypt_Top_sbox_and_1_cse_8_sva_1
      ^ state_4_3_63_32_sva_18 ^ xor_cse_1555 ^ xor_cse_1556 ^ Encrypt_Top_sbox_and_1_cse_50_sva_1
      ^ xor_cse_990 ^ xor_cse_1558 ^ xor_cse_1559;
  assign xor_cse_1562 = plaintext_31_0_sva_16 ^ state_3_3_31_0_sva_16 ^ state_4_3_31_0_sva_16
      ^ state_2_16_1_lpi_4;
  assign xor_cse_1565 = state_2_16_1_lpi_4 & state_3_3_31_0_sva_16;
  assign xor_cse_1566 = state_3_3_31_0_sva_16 & plaintext_31_0_sva_16;
  assign xor_cse_1564 = xor_cse_1565 ^ xor_cse_1566 ^ Encrypt_Top_sbox_and_1_cse_16_sva_1
      ^ state_0_16_lpi_6;
  assign xor_cse_1568 = state_2_58_1_lpi_4 & state_3_3_63_32_sva_26;
  assign xor_cse_1569 = state_3_3_63_32_sva_26 & plaintext_63_32_sva_26;
  assign xor_cse_1567 = state_4_3_63_32_sva_26 ^ xor_cse_1568 ^ xor_cse_1569 ^ Encrypt_Top_sbox_and_1_cse_58_sva_1;
  assign state_1_1_31_0_sva_1_19_1 = xor_cse_1059 ^ xor_cse_1517 ^ xor_cse_1562 ^
      xor_cse_1513 ^ xor_cse_1564 ^ xor_cse_1567;
  assign xor_cse_1571 = state_2_51_1_lpi_4 & state_3_3_63_32_sva_19;
  assign xor_cse_1572 = state_3_3_63_32_sva_19 & plaintext_63_32_sva_19;
  assign xor_cse_1574 = plaintext_31_0_sva_12 ^ state_3_3_31_0_sva_12 ^ state_4_3_31_0_sva_12
      ^ state_2_12_1_lpi_4;
  assign xor_cse_1576 = state_2_12_1_lpi_4 & state_3_3_31_0_sva_12;
  assign xor_cse_1577 = state_3_3_31_0_sva_12 & plaintext_31_0_sva_12;
  assign xor_cse_1575 = xor_cse_1576 ^ xor_cse_1577 ^ Encrypt_Top_sbox_and_1_cse_12_sva_1
      ^ state_0_12_lpi_6;
  assign state_1_1_31_0_sva_1_12_1 = xor_cse_1519 ^ Encrypt_Top_sbox_and_1_cse_9_sva_1
      ^ state_4_3_63_32_sva_19 ^ xor_cse_1571 ^ xor_cse_1572 ^ Encrypt_Top_sbox_and_1_cse_51_sva_1
      ^ xor_cse_1000 ^ xor_cse_1574 ^ xor_cse_1575;
  assign xor_cse_1578 = plaintext_31_0_sva_15 ^ state_3_3_31_0_sva_15 ^ state_4_3_31_0_sva_15
      ^ state_2_15_1_lpi_4;
  assign xor_cse_1581 = state_2_15_1_lpi_4 & state_3_3_31_0_sva_15;
  assign xor_cse_1582 = state_3_3_31_0_sva_15 & plaintext_31_0_sva_15;
  assign xor_cse_1580 = xor_cse_1581 ^ xor_cse_1582 ^ Encrypt_Top_sbox_and_1_cse_15_sva_1
      ^ state_0_15_lpi_6;
  assign xor_cse_1584 = state_2_57_1_lpi_4 & state_3_3_63_32_sva_25;
  assign xor_cse_1585 = state_3_3_63_32_sva_25 & plaintext_63_32_sva_25;
  assign xor_cse_1583 = state_4_3_63_32_sva_25 ^ xor_cse_1584 ^ xor_cse_1585 ^ Encrypt_Top_sbox_and_1_cse_57_sva_1;
  assign state_1_1_31_0_sva_1_18_1 = xor_cse_1050 ^ xor_cse_1535 ^ xor_cse_1578 ^
      xor_cse_1531 ^ xor_cse_1580 ^ xor_cse_1583;
  assign xor_cse_1586 = plaintext_31_0_sva_13 ^ state_3_3_31_0_sva_13 ^ state_4_3_31_0_sva_13
      ^ state_2_13_1_lpi_4;
  assign xor_cse_1588 = state_2_13_1_lpi_4 & state_3_3_31_0_sva_13;
  assign xor_cse_1589 = state_3_3_31_0_sva_13 & plaintext_31_0_sva_13;
  assign xor_cse_1587 = xor_cse_1588 ^ xor_cse_1589 ^ Encrypt_Top_sbox_and_1_cse_13_sva_1
      ^ state_0_13_lpi_6;
  assign xor_cse_1591 = state_4_3_63_32_sva_20 ^ (state_2_52_1_lpi_4 & state_3_3_63_32_sva_20)
      ^ (state_3_3_63_32_sva_20 & plaintext_63_32_sva_20) ^ Encrypt_Top_sbox_and_1_cse_52_sva_1;
  assign state_1_1_31_0_sva_1_13_1 = xor_cse_1009 ^ xor_cse_1540 ^ xor_cse_1586 ^
      xor_cse_1587 ^ xor_cse_1541 ^ xor_cse_1591;
  assign xor_cse_1595 = state_2_56_1_lpi_4 & state_3_3_63_32_sva_24;
  assign xor_cse_1596 = state_3_3_63_32_sva_24 & plaintext_63_32_sva_24;
  assign xor_cse_1598 = plaintext_31_0_sva_14 ^ state_3_3_31_0_sva_14 ^ state_4_3_31_0_sva_14
      ^ state_2_14_1_lpi_4;
  assign xor_cse_1600 = state_2_14_1_lpi_4 & state_3_3_31_0_sva_14;
  assign xor_cse_1601 = state_3_3_31_0_sva_14 & plaintext_31_0_sva_14;
  assign state_1_1_31_0_sva_1_17_1 = xor_cse_1546 ^ state_0_14_lpi_6 ^ state_4_3_63_32_sva_24
      ^ xor_cse_1595 ^ xor_cse_1596 ^ Encrypt_Top_sbox_and_1_cse_56_sva_1 ^ xor_cse_1041
      ^ xor_cse_1598 ^ Encrypt_Top_sbox_and_1_cse_17_sva_1 ^ xor_cse_1600 ^ xor_cse_1601
      ^ Encrypt_Top_sbox_and_1_cse_14_sva_1;
  assign xor_cse_1602 = xor_cse_1600 ^ xor_cse_1601 ^ Encrypt_Top_sbox_and_1_cse_14_sva_1
      ^ state_0_14_lpi_6;
  assign xor_cse_1604 = state_4_3_63_32_sva_21 ^ (state_2_53_1_lpi_4 & state_3_3_63_32_sva_21)
      ^ (state_3_3_63_32_sva_21 & plaintext_63_32_sva_21) ^ Encrypt_Top_sbox_and_1_cse_53_sva_1;
  assign state_1_1_31_0_sva_1_14_1 = xor_cse_1016 ^ xor_cse_1558 ^ xor_cse_1598 ^
      xor_cse_1602 ^ xor_cse_1559 ^ xor_cse_1604;
  assign xor_cse_1609 = state_4_3_63_32_sva_23 ^ (state_2_55_1_lpi_4 & state_3_3_63_32_sva_23)
      ^ (state_3_3_63_32_sva_23 & plaintext_63_32_sva_23) ^ Encrypt_Top_sbox_and_1_cse_55_sva_1;
  assign state_1_1_31_0_sva_1_16_1 = xor_cse_1030 ^ xor_cse_1586 ^ xor_cse_1562 ^
      xor_cse_1564 ^ xor_cse_1587 ^ xor_cse_1609;
  assign xor_cse_1614 = state_4_3_63_32_sva_22 ^ (state_2_54_1_lpi_4 & state_3_3_63_32_sva_22)
      ^ (state_3_3_63_32_sva_22 & plaintext_63_32_sva_22) ^ Encrypt_Top_sbox_and_1_cse_54_sva_1;
  assign state_1_1_31_0_sva_1_15_1 = xor_cse_1021 ^ xor_cse_1574 ^ xor_cse_1578 ^
      xor_cse_1580 ^ xor_cse_1575 ^ xor_cse_1614;
  assign xor_cse_1617 = xor_cse_859 ^ state_4_3_63_32_sva_6 ^ (state_2_38_1_lpi_4
      & state_3_3_63_32_sva_6) ^ (state_3_3_63_32_sva_6 & plaintext_63_32_sva_6);
  assign state_1_1_63_32_sva_1_31_1 = xor_cse_1527 ^ xor_cse_1617 ^ xor_cse_1103
      ^ xor_cse_1490 ^ Encrypt_Top_sbox_and_1_cse_60_sva_1 ^ Encrypt_Top_sbox_and_1_cse_38_sva_1;
  assign xor_cse_1623 = xor_cse_401 ^ state_4_3_63_32_sva_0 ^ (state_2_32_1_lpi_4
      & state_3_3_63_32_sva_0) ^ (state_3_3_63_32_sva_0 & plaintext_63_32_sva_0);
  assign state_1_1_63_32_sva_1_0_1 = xor_cse_1491 ^ xor_cse_1623 ^ xor_cse_1415 ^
      Encrypt_Top_sbox_and_1_cse_32_sva_1 ^ xor_cse_1418 ^ xor_cse_1419 ^ Encrypt_Top_sbox_and_1_cse_29_sva_1
      ^ state_0_29_lpi_6 ^ xor_cse_1497 ^ xor_cse_1498;
  assign xor_cse_1629 = xor_cse_950 ^ state_4_3_63_32_sva_5 ^ (state_2_37_1_lpi_4
      & state_3_3_63_32_sva_5) ^ (state_3_3_63_32_sva_5 & plaintext_63_32_sva_5);
  assign state_1_1_63_32_sva_1_30_1 = xor_cse_1629 ^ xor_cse_1399 ^ xor_cse_1068
      ^ Encrypt_Top_sbox_and_1_cse_62_sva_1 ^ state_4_3_63_32_sva_27 ^ xor_cse_1550
      ^ xor_cse_1551 ^ Encrypt_Top_sbox_and_1_cse_59_sva_1 ^ Encrypt_Top_sbox_and_1_cse_37_sva_1;
  assign xor_cse_1637 = state_4_3_63_32_sva_1 ^ (state_2_33_1_lpi_4 & state_3_3_63_32_sva_1)
      ^ (state_3_3_63_32_sva_1 & plaintext_63_32_sva_1) ^ Encrypt_Top_sbox_and_1_cse_33_sva_1;
  assign state_1_1_63_32_sva_1_1_1 = xor_cse_1505 ^ xor_cse_1393 ^ Encrypt_Top_sbox_and_1_cse_8_sva_1
      ^ xor_cse_419 ^ xor_cse_1391 ^ xor_cse_1637;
  assign xor_cse_1641 = state_2_36_1_lpi_4 & state_3_3_63_32_sva_4;
  assign xor_cse_1642 = state_3_3_63_32_sva_4 & plaintext_63_32_sva_4;
  assign state_1_1_63_32_sva_1_29_1 = xor_cse_1374 ^ Encrypt_Top_sbox_and_1_cse_58_sva_1
      ^ state_4_3_63_32_sva_4 ^ xor_cse_1641 ^ xor_cse_1642 ^ Encrypt_Top_sbox_and_1_cse_36_sva_1
      ^ xor_cse_1059 ^ xor_cse_936 ^ Encrypt_Top_sbox_and_1_cse_61_sva_1 ^ state_4_3_63_32_sva_26
      ^ xor_cse_1568 ^ xor_cse_1569;
  assign xor_cse_1648 = state_2_34_1_lpi_4 & state_3_3_63_32_sva_2;
  assign xor_cse_1649 = state_3_3_63_32_sva_2 & plaintext_63_32_sva_2;
  assign xor_cse_1647 = state_4_3_63_32_sva_2 ^ xor_cse_1648 ^ xor_cse_1649 ^ Encrypt_Top_sbox_and_1_cse_34_sva_1;
  assign state_1_1_63_32_sva_1_2_1 = xor_cse_1519 ^ xor_cse_1368 ^ Encrypt_Top_sbox_and_1_cse_9_sva_1
      ^ xor_cse_431 ^ xor_cse_1367 ^ xor_cse_1647;
  assign xor_cse_1650 = xor_cse_446 ^ state_4_3_63_32_sva_3 ^ (state_2_35_1_lpi_4
      & state_3_3_63_32_sva_3) ^ (state_3_3_63_32_sva_3 & plaintext_63_32_sva_3);
  assign state_1_1_63_32_sva_1_28_1 = xor_cse_1527 ^ xor_cse_1650 ^ xor_cse_1050
      ^ Encrypt_Top_sbox_and_1_cse_60_sva_1 ^ state_4_3_63_32_sva_25 ^ xor_cse_1584
      ^ xor_cse_1585 ^ Encrypt_Top_sbox_and_1_cse_57_sva_1 ^ Encrypt_Top_sbox_and_1_cse_35_sva_1;
  assign state_1_1_63_32_sva_1_3_1 = xor_cse_1623 ^ xor_cse_1650 ^ xor_cse_1540 ^
      Encrypt_Top_sbox_and_1_cse_35_sva_1 ^ Encrypt_Top_sbox_and_1_cse_32_sva_1 ^
      xor_cse_1542 ^ xor_cse_1543 ^ Encrypt_Top_sbox_and_1_cse_10_sva_1 ^ state_0_10_lpi_6;
  assign xor_cse_1660 = state_4_3_63_32_sva_24 ^ xor_cse_1595 ^ xor_cse_1596 ^ Encrypt_Top_sbox_and_1_cse_56_sva_1;
  assign state_1_1_63_32_sva_1_27_1 = xor_cse_1068 ^ xor_cse_1041 ^ xor_cse_431 ^
      state_4_3_63_32_sva_27 ^ xor_cse_1550 ^ xor_cse_1551 ^ Encrypt_Top_sbox_and_1_cse_59_sva_1
      ^ xor_cse_1660 ^ xor_cse_1647;
  assign xor_cse_1662 = state_4_3_63_32_sva_4 ^ xor_cse_1641 ^ xor_cse_1642 ^ Encrypt_Top_sbox_and_1_cse_36_sva_1;
  assign state_1_1_63_32_sva_1_4_1 = xor_cse_936 ^ xor_cse_419 ^ xor_cse_1558 ^ xor_cse_1662
      ^ xor_cse_1637 ^ xor_cse_1559;
  assign state_1_1_63_32_sva_1_26_1 = xor_cse_1059 ^ xor_cse_1030 ^ xor_cse_419 ^
      xor_cse_1567 ^ xor_cse_1609 ^ xor_cse_1637;
  assign state_1_1_63_32_sva_1_5_1 = xor_cse_1629 ^ Encrypt_Top_sbox_and_1_cse_34_sva_1
      ^ xor_cse_1576 ^ xor_cse_1577 ^ Encrypt_Top_sbox_and_1_cse_12_sva_1 ^ state_0_12_lpi_6
      ^ xor_cse_431 ^ xor_cse_1574 ^ Encrypt_Top_sbox_and_1_cse_37_sva_1 ^ state_4_3_63_32_sva_2
      ^ xor_cse_1648 ^ xor_cse_1649;
  assign state_1_1_63_32_sva_1_25_1 = xor_cse_1623 ^ xor_cse_1614 ^ Encrypt_Top_sbox_and_1_cse_32_sva_1
      ^ xor_cse_1050 ^ xor_cse_1021 ^ xor_cse_1583;
  assign state_1_1_63_32_sva_1_6_1 = xor_cse_1617 ^ xor_cse_1650 ^ xor_cse_1586 ^
      Encrypt_Top_sbox_and_1_cse_38_sva_1 ^ Encrypt_Top_sbox_and_1_cse_35_sva_1 ^
      xor_cse_1588 ^ xor_cse_1589 ^ Encrypt_Top_sbox_and_1_cse_13_sva_1 ^ state_0_13_lpi_6;
  assign state_1_1_63_32_sva_1_24_1 = xor_cse_1041 ^ xor_cse_1016 ^ xor_cse_1367
      ^ xor_cse_1660 ^ xor_cse_1604 ^ xor_cse_1368;
  assign xor_cse_1680 = state_4_3_63_32_sva_7 ^ xor_cse_1384 ^ xor_cse_1385 ^ Encrypt_Top_sbox_and_1_cse_39_sva_1;
  assign state_1_1_63_32_sva_1_7_1 = xor_cse_936 ^ xor_cse_867 ^ xor_cse_1598 ^ xor_cse_1680
      ^ xor_cse_1662 ^ xor_cse_1602;
  assign state_1_1_63_32_sva_1_23_1 = xor_cse_1030 ^ xor_cse_1009 ^ xor_cse_1391
      ^ xor_cse_1609 ^ xor_cse_1591 ^ xor_cse_1393;
  assign state_1_1_63_32_sva_1_8_1 = xor_cse_1629 ^ xor_cse_1403 ^ xor_cse_1578 ^
      Encrypt_Top_sbox_and_1_cse_40_sva_1 ^ Encrypt_Top_sbox_and_1_cse_37_sva_1 ^
      xor_cse_1581 ^ xor_cse_1582 ^ Encrypt_Top_sbox_and_1_cse_15_sva_1 ^ state_0_15_lpi_6;
  assign xor_cse_1690 = state_4_3_63_32_sva_19 ^ xor_cse_1571 ^ xor_cse_1572 ^ Encrypt_Top_sbox_and_1_cse_51_sva_1;
  assign state_1_1_63_32_sva_1_22_1 = xor_cse_1000 ^ xor_cse_1021 ^ xor_cse_1415
      ^ xor_cse_1614 ^ xor_cse_1690 ^ xor_cse_1417;
  assign state_1_1_63_32_sva_1_9_1 = xor_cse_1617 ^ xor_cse_1423 ^ xor_cse_1562 ^
      Encrypt_Top_sbox_and_1_cse_41_sva_1 ^ Encrypt_Top_sbox_and_1_cse_38_sva_1 ^
      xor_cse_1565 ^ xor_cse_1566 ^ Encrypt_Top_sbox_and_1_cse_16_sva_1 ^ state_0_16_lpi_6;
  assign xor_cse_1696 = state_4_3_63_32_sva_18 ^ xor_cse_1555 ^ xor_cse_1556 ^ Encrypt_Top_sbox_and_1_cse_50_sva_1;
  assign state_1_1_63_32_sva_1_21_1 = xor_cse_990 ^ xor_cse_1016 ^ xor_cse_1366 ^
      xor_cse_1604 ^ xor_cse_1696 ^ xor_cse_1371;
  assign state_1_1_63_32_sva_1_10_1 = xor_cse_1546 ^ xor_cse_1680 ^ Encrypt_Top_sbox_and_1_cse_17_sva_1
      ^ xor_cse_899 ^ xor_cse_867 ^ xor_cse_1446;
  assign xor_cse_1702 = state_4_3_63_32_sva_17 ^ xor_cse_1545 ^ xor_cse_1538 ^ Encrypt_Top_sbox_and_1_cse_49_sva_1;
  assign state_1_1_63_32_sva_1_20_1 = xor_cse_1009 ^ xor_cse_981 ^ xor_cse_1392 ^
      xor_cse_1591 ^ xor_cse_1702 ^ xor_cse_1396;
  assign state_1_1_63_32_sva_1_11_1 = xor_cse_1456 ^ xor_cse_1403 ^ xor_cse_1535
      ^ Encrypt_Top_sbox_and_1_cse_43_sva_1 ^ Encrypt_Top_sbox_and_1_cse_40_sva_1
      ^ xor_cse_1532 ^ xor_cse_1533 ^ Encrypt_Top_sbox_and_1_cse_18_sva_1 ^ state_0_18_lpi_6;
  assign xor_cse_1708 = state_4_3_63_32_sva_16 ^ xor_cse_1525 ^ xor_cse_1526 ^ Encrypt_Top_sbox_and_1_cse_48_sva_1;
  assign state_1_1_63_32_sva_1_19_1 = xor_cse_1000 ^ xor_cse_970 ^ xor_cse_1416 ^
      xor_cse_1690 ^ xor_cse_1708 ^ xor_cse_1420;
  assign state_1_1_63_32_sva_1_12_1 = xor_cse_1468 ^ xor_cse_1423 ^ xor_cse_1517
      ^ Encrypt_Top_sbox_and_1_cse_44_sva_1 ^ Encrypt_Top_sbox_and_1_cse_41_sva_1
      ^ xor_cse_1514 ^ xor_cse_1515 ^ Encrypt_Top_sbox_and_1_cse_19_sva_1 ^ state_0_19_lpi_6;
  assign xor_cse_1714 = state_4_3_63_32_sva_15 ^ xor_cse_1511 ^ xor_cse_1512 ^ Encrypt_Top_sbox_and_1_cse_47_sva_1;
  assign state_1_1_63_32_sva_1_18_1 = xor_cse_990 ^ xor_cse_961 ^ xor_cse_1439 ^
      xor_cse_1696 ^ xor_cse_1714 ^ xor_cse_1441;
  assign state_1_1_63_32_sva_1_13_1 = xor_cse_899 ^ xor_cse_935 ^ xor_cse_1503 ^
      xor_cse_1482 ^ xor_cse_1446 ^ xor_cse_1499;
  assign state_1_1_63_32_sva_1_17_1 = xor_cse_1492 ^ Encrypt_Top_sbox_and_1_cse_46_sva_1
      ^ xor_cse_1454 ^ xor_cse_1455 ^ Encrypt_Top_sbox_and_1_cse_24_sva_1 ^ state_0_24_lpi_6
      ^ xor_cse_981 ^ xor_cse_1451 ^ xor_cse_1702;
  assign state_1_1_63_32_sva_1_14_1 = xor_cse_1456 ^ xor_cse_1492 ^ xor_cse_1485
      ^ Encrypt_Top_sbox_and_1_cse_46_sva_1 ^ Encrypt_Top_sbox_and_1_cse_43_sva_1
      ^ xor_cse_1488 ^ xor_cse_1489 ^ Encrypt_Top_sbox_and_1_cse_21_sva_1 ^ state_0_21_lpi_6;
  assign state_1_1_63_32_sva_1_16_1 = xor_cse_935 ^ xor_cse_970 ^ xor_cse_1463 ^
      xor_cse_1708 ^ xor_cse_1482 ^ xor_cse_1465;
  assign state_1_1_63_32_sva_1_15_1 = xor_cse_1468 ^ Encrypt_Top_sbox_and_1_cse_44_sva_1
      ^ xor_cse_1478 ^ xor_cse_1479 ^ Encrypt_Top_sbox_and_1_cse_22_sva_1 ^ state_0_22_lpi_6
      ^ xor_cse_961 ^ xor_cse_1475 ^ xor_cse_1714;
  assign xor_cse_1731 = state_4_3_63_32_sva_8 ^ plaintext_63_32_sva_8 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_8
      ^ state_3_3_63_32_sva_8;
  assign xor_cse_1732 = state_4_3_63_32_sva_31 ^ plaintext_63_32_sva_31 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_31
      ^ state_3_3_63_32_sva_31;
  assign xor_cse_1734 = plaintext_31_0_sva_6 ^ state_4_3_31_0_sva_6 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_6
      ^ state_3_3_31_0_sva_6;
  assign xor_cse_1733 = Encrypt_Top_sbox_and_2_cse_6_sva_1 ^ xor_cse_1734 ^ Encrypt_Top_sbox_and_2_cse_63_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_40_sva_1;
  assign xor_cse_1735 = plaintext_31_0_sva_7 ^ state_4_3_31_0_sva_7 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_7
      ^ state_3_3_31_0_sva_7;
  assign xor_cse_1736 = state_4_3_63_32_sva_9 ^ plaintext_63_32_sva_9 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_9
      ^ state_3_3_63_32_sva_9;
  assign xor_cse_1738 = plaintext_31_0_sva_0 ^ state_4_3_31_0_sva_0 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_0
      ^ state_3_3_31_0_sva_0;
  assign xor_cse_1737 = Encrypt_Top_sbox_and_2_cse_0_sva_1 ^ xor_cse_1738 ^ Encrypt_Top_sbox_and_2_cse_7_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_41_sva_1;
  assign xor_cse_1739 = state_4_3_63_32_sva_7 ^ plaintext_63_32_sva_7 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_7
      ^ state_3_3_63_32_sva_7;
  assign xor_cse_1741 = plaintext_31_0_sva_5 ^ state_4_3_31_0_sva_5 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_5
      ^ state_3_3_31_0_sva_5;
  assign xor_cse_1740 = Encrypt_Top_sbox_and_2_cse_5_sva_1 ^ xor_cse_1741 ^ state_4_3_63_32_sva_30
      ^ Encrypt_Top_sbox_and_2_cse_39_sva_1;
  assign xor_cse_1742 = state_4_3_63_32_sva_10 ^ plaintext_63_32_sva_10 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_10
      ^ state_3_3_63_32_sva_10;
  assign xor_cse_1743 = state_4_3_31_0_sva_8 ^ plaintext_31_0_sva_8 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_8
      ^ state_3_3_31_0_sva_8;
  assign xor_cse_1745 = plaintext_31_0_sva_1 ^ state_4_3_31_0_sva_1 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_1
      ^ state_3_3_31_0_sva_1;
  assign xor_cse_1744 = Encrypt_Top_sbox_and_2_cse_1_sva_1 ^ xor_cse_1745 ^ Encrypt_Top_sbox_and_2_cse_8_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_42_sva_1;
  assign xor_cse_1746 = state_4_3_63_32_sva_6 ^ plaintext_63_32_sva_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_6
      ^ state_3_3_63_32_sva_6;
  assign xor_cse_1748 = plaintext_31_0_sva_4 ^ state_4_3_31_0_sva_4 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_4
      ^ state_3_3_31_0_sva_4;
  assign xor_cse_1747 = Encrypt_Top_sbox_and_2_cse_4_sva_1 ^ xor_cse_1748 ^ state_4_3_63_32_sva_29
      ^ Encrypt_Top_sbox_and_2_cse_38_sva_1;
  assign xor_cse_1749 = state_4_3_63_32_sva_11 ^ plaintext_63_32_sva_11 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_11
      ^ state_3_3_63_32_sva_11;
  assign xor_cse_1750 = state_4_3_31_0_sva_9 ^ plaintext_31_0_sva_9 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_9
      ^ state_3_3_31_0_sva_9;
  assign xor_cse_1752 = plaintext_31_0_sva_2 ^ state_4_3_31_0_sva_2 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_2
      ^ state_3_3_31_0_sva_2;
  assign xor_cse_1751 = Encrypt_Top_sbox_and_2_cse_2_sva_1 ^ xor_cse_1752 ^ Encrypt_Top_sbox_and_2_cse_9_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_43_sva_1;
  assign xor_cse_1753 = state_4_3_63_32_sva_5 ^ plaintext_63_32_sva_5 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_5
      ^ state_3_3_63_32_sva_5;
  assign xor_cse_1755 = plaintext_31_0_sva_3 ^ state_4_3_31_0_sva_3 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_3
      ^ state_3_3_31_0_sva_3;
  assign xor_cse_1754 = Encrypt_Top_sbox_and_2_cse_3_sva_1 ^ xor_cse_1755 ^ state_4_3_63_32_sva_28
      ^ Encrypt_Top_sbox_and_2_cse_37_sva_1;
  assign xor_cse_1756 = state_4_3_63_32_sva_12 ^ plaintext_63_32_sva_12 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_12
      ^ state_3_3_63_32_sva_12;
  assign xor_cse_1757 = state_4_3_31_0_sva_10 ^ xor_cse_861 ^ Encrypt_Top_sbox_and_2_cse_3_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_44_sva_1;
  assign xor_cse_1758 = state_4_3_63_32_sva_27 ^ plaintext_63_32_sva_27 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_27
      ^ state_3_3_63_32_sva_27;
  assign xor_cse_1760 = state_4_3_63_32_sva_4 ^ plaintext_63_32_sva_4 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_4
      ^ state_3_3_63_32_sva_4;
  assign xor_cse_1759 = Encrypt_Top_sbox_and_2_cse_36_sva_1 ^ xor_cse_1760 ^ Encrypt_Top_sbox_and_2_cse_59_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_2_sva_1;
  assign xor_cse_1761 = state_4_3_63_32_sva_13 ^ plaintext_63_32_sva_13 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_13
      ^ state_3_3_63_32_sva_13;
  assign xor_cse_1762 = state_4_3_31_0_sva_11 ^ xor_cse_868 ^ Encrypt_Top_sbox_and_2_cse_4_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_45_sva_1;
  assign xor_cse_1763 = state_4_3_63_32_sva_26 ^ plaintext_63_32_sva_26 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_26
      ^ state_3_3_63_32_sva_26;
  assign xor_cse_1765 = state_4_3_63_32_sva_3 ^ plaintext_63_32_sva_3 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_3
      ^ state_3_3_63_32_sva_3;
  assign xor_cse_1764 = Encrypt_Top_sbox_and_2_cse_35_sva_1 ^ xor_cse_1765 ^ Encrypt_Top_sbox_and_2_cse_58_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_1_sva_1;
  assign xor_cse_1766 = state_4_3_63_32_sva_14 ^ plaintext_63_32_sva_14 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_14
      ^ state_3_3_63_32_sva_14;
  assign xor_cse_1767 = state_4_3_31_0_sva_12 ^ xor_cse_880 ^ Encrypt_Top_sbox_and_2_cse_5_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_46_sva_1;
  assign xor_cse_1768 = state_4_3_63_32_sva_25 ^ plaintext_63_32_sva_25 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_25
      ^ state_3_3_63_32_sva_25;
  assign xor_cse_1770 = state_4_3_63_32_sva_2 ^ plaintext_63_32_sva_2 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_2
      ^ state_3_3_63_32_sva_2;
  assign xor_cse_1769 = Encrypt_Top_sbox_and_2_cse_34_sva_1 ^ xor_cse_1770 ^ Encrypt_Top_sbox_and_2_cse_57_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_0_sva_1;
  assign xor_cse_1771 = state_4_3_63_32_sva_15 ^ plaintext_63_32_sva_15 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_15
      ^ state_3_3_63_32_sva_15;
  assign xor_cse_1772 = state_4_3_31_0_sva_13 ^ xor_cse_890 ^ Encrypt_Top_sbox_and_2_cse_6_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_47_sva_1;
  assign xor_cse_1773 = state_4_3_63_32_sva_24 ^ plaintext_63_32_sva_24 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_24
      ^ state_3_3_63_32_sva_24;
  assign xor_cse_1775 = state_4_3_63_32_sva_1 ^ plaintext_63_32_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_1
      ^ state_3_3_63_32_sva_1;
  assign xor_cse_1774 = Encrypt_Top_sbox_and_2_cse_33_sva_1 ^ xor_cse_1775 ^ Encrypt_Top_sbox_and_2_cse_56_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_63_sva_1;
  assign xor_cse_1776 = state_4_3_63_32_sva_16 ^ plaintext_63_32_sva_16 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_16
      ^ state_3_3_63_32_sva_16;
  assign xor_cse_1777 = state_4_3_31_0_sva_14 ^ xor_cse_900 ^ Encrypt_Top_sbox_and_2_cse_7_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_48_sva_1;
  assign xor_cse_1778 = state_4_3_63_32_sva_23 ^ plaintext_63_32_sva_23 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_23
      ^ state_3_3_63_32_sva_23;
  assign xor_cse_1780 = state_4_3_63_32_sva_0 ^ plaintext_63_32_sva_0 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_0
      ^ state_3_3_63_32_sva_0;
  assign xor_cse_1779 = Encrypt_Top_sbox_and_2_cse_32_sva_1 ^ xor_cse_1780 ^ Encrypt_Top_sbox_and_2_cse_55_sva_1
      ^ state_4_3_63_32_sva_30;
  assign xor_cse_1781 = state_4_3_63_32_sva_17 ^ plaintext_63_32_sva_17 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_17
      ^ state_3_3_63_32_sva_17;
  assign xor_cse_1782 = state_4_3_31_0_sva_15 ^ xor_cse_912 ^ Encrypt_Top_sbox_and_2_cse_8_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_49_sva_1;
  assign xor_cse_1783 = state_4_3_63_32_sva_22 ^ plaintext_63_32_sva_22 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_22
      ^ state_3_3_63_32_sva_22;
  assign xor_cse_1784 = state_4_3_31_0_sva_31 ^ xor_cse_390 ^ Encrypt_Top_sbox_and_2_cse_54_sva_1
      ^ state_4_3_63_32_sva_29;
  assign xor_cse_1785 = state_4_3_63_32_sva_18 ^ plaintext_63_32_sva_18 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_18
      ^ state_3_3_63_32_sva_18;
  assign xor_cse_1786 = state_4_3_31_0_sva_16 ^ xor_cse_926 ^ Encrypt_Top_sbox_and_2_cse_9_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_50_sva_1;
  assign xor_cse_1787 = state_4_3_63_32_sva_21 ^ plaintext_63_32_sva_21 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_21
      ^ state_3_3_63_32_sva_21;
  assign xor_cse_1788 = state_4_3_31_0_sva_30 ^ xor_cse_379 ^ Encrypt_Top_sbox_and_2_cse_53_sva_1
      ^ state_4_3_63_32_sva_28;
  assign xor_cse_1789 = state_4_3_63_32_sva_19 ^ plaintext_63_32_sva_19 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_19
      ^ state_3_3_63_32_sva_19;
  assign xor_cse_1790 = state_4_3_31_0_sva_17 ^ plaintext_31_0_sva_17 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_17
      ^ state_3_3_31_0_sva_17;
  assign xor_cse_1792 = state_4_3_63_32_sva_20 ^ plaintext_63_32_sva_20 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_20
      ^ state_3_3_63_32_sva_20;
  assign xor_cse_1793 = state_4_3_31_0_sva_29 ^ xor_cse_366 ^ Encrypt_Top_sbox_and_2_cse_52_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_59_sva_1;
  assign xor_cse_1794 = state_4_3_31_0_sva_18 ^ xor_cse_951 ^ state_4_3_31_0_sva_11
      ^ Encrypt_Top_sbox_and_2_cse_52_sva_1;
  assign xor_cse_1795 = state_4_3_31_0_sva_28 ^ xor_cse_354 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_58_sva_1;
  assign xor_cse_1796 = state_4_3_31_0_sva_19 ^ xor_cse_350 ^ state_4_3_31_0_sva_12
      ^ Encrypt_Top_sbox_and_2_cse_53_sva_1;
  assign xor_cse_1797 = state_4_3_31_0_sva_27 ^ xor_cse_1031 ^ Encrypt_Top_sbox_and_2_cse_50_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_57_sva_1;
  assign xor_cse_1798 = state_4_3_31_0_sva_20 ^ xor_cse_362 ^ state_4_3_31_0_sva_13
      ^ Encrypt_Top_sbox_and_2_cse_54_sva_1;
  assign xor_cse_1799 = state_4_3_31_0_sva_26 ^ xor_cse_448 ^ Encrypt_Top_sbox_and_2_cse_49_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_56_sva_1;
  assign xor_cse_1800 = state_4_3_31_0_sva_21 ^ xor_cse_375 ^ state_4_3_31_0_sva_14
      ^ Encrypt_Top_sbox_and_2_cse_55_sva_1;
  assign xor_cse_1801 = state_4_3_31_0_sva_25 ^ xor_cse_428 ^ Encrypt_Top_sbox_and_2_cse_48_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_55_sva_1;
  assign xor_cse_1802 = state_4_3_31_0_sva_22 ^ xor_cse_387 ^ state_4_3_31_0_sva_15
      ^ Encrypt_Top_sbox_and_2_cse_56_sva_1;
  assign xor_cse_1803 = state_4_3_31_0_sva_24 ^ xor_cse_415 ^ Encrypt_Top_sbox_and_2_cse_47_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_54_sva_1;
  assign xor_cse_1804 = state_4_3_31_0_sva_23 ^ xor_cse_403 ^ state_4_3_31_0_sva_16
      ^ Encrypt_Top_sbox_and_2_cse_57_sva_1;
  assign xor_cse_1835 = state_0_16_lpi_6 ^ xor_cse_1562 ^ (state_4_3_31_0_sva_16
      & state_0_16_lpi_6) ^ (state_3_3_31_0_sva_16 & state_0_16_lpi_6);
  assign xor_cse_1838 = xor_cse_1103 ^ state_4_3_63_32_sva_31 ^ (state_4_3_63_32_sva_31
      & state_0_63_lpi_6) ^ (state_3_3_63_32_sva_31 & state_0_63_lpi_6);
  assign xor_cse_1843 = state_4_3_31_0_sva_9 & state_0_9_lpi_6;
  assign xor_cse_1844 = state_3_3_31_0_sva_9 & state_0_9_lpi_6;
  assign xor_cse_1842 = xor_cse_1843 ^ xor_cse_1844 ^ state_4_3_31_0_sva_9;
  assign xor_cse_1845 = state_0_10_lpi_6 ^ xor_cse_1540 ^ (state_4_3_31_0_sva_10
      & state_0_10_lpi_6) ^ (state_3_3_31_0_sva_10 & state_0_10_lpi_6);
  assign xor_cse_1849 = plaintext_31_0_sva_0 ^ state_4_3_31_0_sva_0 ^ (state_4_3_31_0_sva_0
      & state_0_0_lpi_6) ^ (state_3_3_31_0_sva_0 & state_0_0_lpi_6);
  assign xor_cse_1853 = state_4_3_31_0_sva_17 & state_0_17_lpi_6;
  assign xor_cse_1854 = state_3_3_31_0_sva_17 & state_0_17_lpi_6;
  assign xor_cse_1852 = xor_cse_1853 ^ xor_cse_1854 ^ state_4_3_31_0_sva_17;
  assign xor_cse_1855 = state_0_15_lpi_6 ^ xor_cse_1578 ^ (state_4_3_31_0_sva_15
      & state_0_15_lpi_6) ^ (state_3_3_31_0_sva_15 & state_0_15_lpi_6);
  assign xor_cse_1860 = state_4_3_63_32_sva_30 & state_0_62_lpi_6;
  assign xor_cse_1861 = state_3_3_63_32_sva_30 & state_0_62_lpi_6;
  assign xor_cse_1862 = state_4_3_31_0_sva_8 & state_0_8_lpi_6;
  assign xor_cse_1859 = state_0_62_lpi_6 ^ xor_cse_1860 ^ xor_cse_1861 ^ xor_cse_1862;
  assign xor_cse_1864 = state_3_3_31_0_sva_8 & state_0_8_lpi_6;
  assign xor_cse_1865 = plaintext_31_0_sva_1 ^ state_4_3_31_0_sva_1 ^ (state_4_3_31_0_sva_1
      & state_0_1_lpi_6) ^ (state_3_3_31_0_sva_1 & state_0_1_lpi_6);
  assign xor_cse_1868 = state_0_11_lpi_6 ^ xor_cse_1558 ^ (state_4_3_31_0_sva_11
      & state_0_11_lpi_6) ^ (state_3_3_31_0_sva_11 & state_0_11_lpi_6);
  assign xor_cse_1871 = state_0_18_lpi_6 ^ xor_cse_1535 ^ (state_4_3_31_0_sva_18
      & state_0_18_lpi_6) ^ (state_3_3_31_0_sva_18 & state_0_18_lpi_6);
  assign xor_cse_1874 = plaintext_31_0_sva_7 ^ state_4_3_31_0_sva_7 ^ (state_4_3_31_0_sva_7
      & state_0_7_lpi_6) ^ (state_3_3_31_0_sva_7 & state_0_7_lpi_6);
  assign xor_cse_1877 = state_0_14_lpi_6 ^ xor_cse_1598 ^ (state_4_3_31_0_sva_14
      & state_0_14_lpi_6) ^ (state_3_3_31_0_sva_14 & state_0_14_lpi_6);
  assign xor_cse_1881 = state_4_3_63_32_sva_29 & state_0_61_lpi_6;
  assign xor_cse_1882 = state_3_3_63_32_sva_29 & state_0_61_lpi_6;
  assign xor_cse_1880 = state_0_61_lpi_6 ^ xor_cse_1881 ^ xor_cse_1882 ^ xor_cse_1375;
  assign xor_cse_1883 = plaintext_31_0_sva_2 ^ state_4_3_31_0_sva_2 ^ (state_4_3_31_0_sva_2
      & state_0_2_lpi_6) ^ (state_3_3_31_0_sva_2 & state_0_2_lpi_6);
  assign xor_cse_1886 = state_0_12_lpi_6 ^ xor_cse_1574 ^ (state_4_3_31_0_sva_12
      & state_0_12_lpi_6) ^ (state_3_3_31_0_sva_12 & state_0_12_lpi_6);
  assign xor_cse_1889 = state_0_19_lpi_6 ^ xor_cse_1517 ^ (state_4_3_31_0_sva_19
      & state_0_19_lpi_6) ^ (state_3_3_31_0_sva_19 & state_0_19_lpi_6);
  assign xor_cse_1892 = plaintext_31_0_sva_6 ^ state_4_3_31_0_sva_6 ^ (state_4_3_31_0_sva_6
      & state_0_6_lpi_6) ^ (state_3_3_31_0_sva_6 & state_0_6_lpi_6);
  assign xor_cse_1895 = state_0_13_lpi_6 ^ xor_cse_1586 ^ (state_4_3_31_0_sva_13
      & state_0_13_lpi_6) ^ (state_3_3_31_0_sva_13 & state_0_13_lpi_6);
  assign xor_cse_1899 = state_4_3_63_32_sva_28 & state_0_60_lpi_6;
  assign xor_cse_1900 = state_3_3_63_32_sva_28 & state_0_60_lpi_6;
  assign xor_cse_1898 = state_0_60_lpi_6 ^ xor_cse_1899 ^ xor_cse_1900 ^ xor_cse_1528;
  assign xor_cse_1901 = plaintext_31_0_sva_3 ^ state_4_3_31_0_sva_3 ^ (state_4_3_31_0_sva_3
      & state_0_3_lpi_6) ^ (state_3_3_31_0_sva_3 & state_0_3_lpi_6);
  assign xor_cse_1904 = state_0_20_lpi_6 ^ xor_cse_1503 ^ (state_4_3_31_0_sva_20
      & state_0_20_lpi_6) ^ (state_3_3_31_0_sva_20 & state_0_20_lpi_6);
  assign xor_cse_1907 = plaintext_31_0_sva_5 ^ state_4_3_31_0_sva_5 ^ (state_4_3_31_0_sva_5
      & state_0_5_lpi_6) ^ (state_3_3_31_0_sva_5 & state_0_5_lpi_6);
  assign xor_cse_1910 = xor_cse_1068 ^ state_4_3_63_32_sva_27 ^ (state_4_3_63_32_sva_27
      & state_0_59_lpi_6) ^ (state_3_3_63_32_sva_27 & state_0_59_lpi_6);
  assign xor_cse_1913 = plaintext_31_0_sva_4 ^ state_4_3_31_0_sva_4 ^ (state_4_3_31_0_sva_4
      & state_0_4_lpi_6) ^ (state_3_3_31_0_sva_4 & state_0_4_lpi_6);
  assign xor_cse_1916 = state_0_21_lpi_6 ^ xor_cse_1485 ^ (state_4_3_31_0_sva_21
      & state_0_21_lpi_6) ^ (state_3_3_31_0_sva_21 & state_0_21_lpi_6);
  assign xor_cse_1919 = xor_cse_1059 ^ state_4_3_63_32_sva_26 ^ (state_4_3_63_32_sva_26
      & state_0_58_lpi_6) ^ (state_3_3_63_32_sva_26 & state_0_58_lpi_6);
  assign xor_cse_1922 = state_0_22_lpi_6 ^ xor_cse_1475 ^ (state_4_3_31_0_sva_22
      & state_0_22_lpi_6) ^ (state_3_3_31_0_sva_22 & state_0_22_lpi_6);
  assign xor_cse_1925 = xor_cse_1050 ^ state_4_3_63_32_sva_25 ^ (state_4_3_63_32_sva_25
      & state_0_57_lpi_6) ^ (state_3_3_63_32_sva_25 & state_0_57_lpi_6);
  assign xor_cse_1928 = state_0_23_lpi_6 ^ xor_cse_1463 ^ (state_4_3_31_0_sva_23
      & state_0_23_lpi_6) ^ (state_3_3_31_0_sva_23 & state_0_23_lpi_6);
  assign xor_cse_1931 = xor_cse_1041 ^ state_4_3_63_32_sva_24 ^ (state_4_3_63_32_sva_24
      & state_0_56_lpi_6) ^ (state_3_3_63_32_sva_24 & state_0_56_lpi_6);
  assign xor_cse_1936 = state_0_24_lpi_6 ^ xor_cse_1451 ^ (state_4_3_31_0_sva_24
      & state_0_24_lpi_6) ^ (state_3_3_31_0_sva_24 & state_0_24_lpi_6);
  assign xor_cse_1941 = xor_cse_1030 ^ state_4_3_63_32_sva_23 ^ (state_4_3_63_32_sva_23
      & state_0_55_lpi_6) ^ (state_3_3_63_32_sva_23 & state_0_55_lpi_6);
  assign xor_cse_1945 = xor_cse_1862 ^ xor_cse_1864 ^ state_4_3_31_0_sva_8;
  assign xor_cse_1946 = state_0_25_lpi_6 ^ xor_cse_1439 ^ (state_4_3_31_0_sva_25
      & state_0_25_lpi_6) ^ (state_3_3_31_0_sva_25 & state_0_25_lpi_6);
  assign xor_cse_1951 = xor_cse_1021 ^ state_4_3_63_32_sva_22 ^ (state_4_3_63_32_sva_22
      & state_0_54_lpi_6) ^ (state_3_3_63_32_sva_22 & state_0_54_lpi_6);
  assign xor_cse_1955 = state_0_26_lpi_6 ^ xor_cse_1416 ^ (state_4_3_31_0_sva_26
      & state_0_26_lpi_6) ^ (state_3_3_31_0_sva_26 & state_0_26_lpi_6);
  assign xor_cse_1960 = xor_cse_1016 ^ state_4_3_63_32_sva_21 ^ (state_4_3_63_32_sva_21
      & state_0_53_lpi_6) ^ (state_3_3_63_32_sva_21 & state_0_53_lpi_6);
  assign xor_cse_1963 = state_0_27_lpi_6 ^ xor_cse_1392 ^ (state_4_3_31_0_sva_27
      & state_0_27_lpi_6) ^ (state_3_3_31_0_sva_27 & state_0_27_lpi_6);
  assign xor_cse_1966 = xor_cse_1009 ^ state_4_3_63_32_sva_20 ^ (state_4_3_63_32_sva_20
      & state_0_52_lpi_6) ^ (state_3_3_63_32_sva_20 & state_0_52_lpi_6);
  assign xor_cse_1969 = state_0_62_lpi_6 ^ xor_cse_1860 ^ xor_cse_1861 ^ xor_cse_1400;
  assign xor_cse_1970 = state_0_28_lpi_6 ^ xor_cse_1366 ^ (state_4_3_31_0_sva_28
      & state_0_28_lpi_6) ^ (state_3_3_31_0_sva_28 & state_0_28_lpi_6);
  assign xor_cse_1973 = xor_cse_1000 ^ state_4_3_63_32_sva_19 ^ (state_4_3_63_32_sva_19
      & state_0_51_lpi_6) ^ (state_3_3_63_32_sva_19 & state_0_51_lpi_6);
  assign xor_cse_1976 = state_0_29_lpi_6 ^ xor_cse_1415 ^ (state_4_3_31_0_sva_29
      & state_0_29_lpi_6) ^ (state_3_3_31_0_sva_29 & state_0_29_lpi_6);
  assign xor_cse_1979 = xor_cse_990 ^ state_4_3_63_32_sva_18 ^ (state_4_3_63_32_sva_18
      & state_0_50_lpi_6) ^ (state_3_3_63_32_sva_18 & state_0_50_lpi_6);
  assign xor_cse_1982 = state_0_30_lpi_6 ^ xor_cse_1391 ^ (state_4_3_31_0_sva_30
      & state_0_30_lpi_6) ^ (state_3_3_31_0_sva_30 & state_0_30_lpi_6);
  assign xor_cse_1985 = xor_cse_981 ^ state_4_3_63_32_sva_17 ^ (state_4_3_63_32_sva_17
      & state_0_49_lpi_6) ^ (state_3_3_63_32_sva_17 & state_0_49_lpi_6);
  assign xor_cse_1988 = state_0_31_lpi_6 ^ xor_cse_1367 ^ (state_4_3_31_0_sva_31
      & state_0_31_lpi_6) ^ (state_3_3_31_0_sva_31 & state_0_31_lpi_6);
  assign xor_cse_1991 = xor_cse_970 ^ state_4_3_63_32_sva_16 ^ (state_4_3_63_32_sva_16
      & state_0_48_lpi_6) ^ (state_3_3_63_32_sva_16 & state_0_48_lpi_6);
  assign xor_cse_1996 = state_4_3_63_32_sva_0 & state_0_32_lpi_6;
  assign xor_cse_1997 = state_3_3_63_32_sva_0 & state_0_32_lpi_6;
  assign xor_cse_1995 = xor_cse_1996 ^ xor_cse_1997 ^ state_4_3_63_32_sva_0;
  assign xor_cse_1998 = xor_cse_961 ^ state_4_3_63_32_sva_15 ^ (state_4_3_63_32_sva_15
      & state_0_47_lpi_6) ^ (state_3_3_63_32_sva_15 & state_0_47_lpi_6);
  assign xor_cse_2001 = xor_cse_419 ^ state_4_3_63_32_sva_1 ^ (state_4_3_63_32_sva_1
      & state_0_33_lpi_6) ^ (state_3_3_63_32_sva_1 & state_0_33_lpi_6);
  assign xor_cse_2006 = state_4_3_63_32_sva_14 & state_0_46_lpi_6;
  assign xor_cse_2007 = state_3_3_63_32_sva_14 & state_0_46_lpi_6;
  assign xor_cse_2005 = xor_cse_2006 ^ xor_cse_2007 ^ state_4_3_63_32_sva_14;
  assign xor_cse_2008 = xor_cse_431 ^ state_4_3_63_32_sva_2 ^ (state_4_3_63_32_sva_2
      & state_0_34_lpi_6) ^ (state_3_3_63_32_sva_2 & state_0_34_lpi_6);
  assign xor_cse_2013 = xor_cse_935 ^ state_4_3_63_32_sva_13 ^ (state_4_3_63_32_sva_13
      & state_0_45_lpi_6) ^ (state_3_3_63_32_sva_13 & state_0_45_lpi_6);
  assign xor_cse_2018 = state_4_3_63_32_sva_3 & state_0_35_lpi_6;
  assign xor_cse_2019 = state_3_3_63_32_sva_3 & state_0_35_lpi_6;
  assign xor_cse_2017 = xor_cse_2018 ^ xor_cse_2019 ^ state_4_3_63_32_sva_3;
  assign xor_cse_2022 = state_4_3_63_32_sva_12 & state_0_44_lpi_6;
  assign xor_cse_2021 = state_0_61_lpi_6 ^ xor_cse_1881 ^ xor_cse_1882 ^ xor_cse_2022;
  assign xor_cse_2024 = state_3_3_63_32_sva_12 & state_0_44_lpi_6;
  assign xor_cse_2025 = xor_cse_936 ^ state_4_3_63_32_sva_4 ^ (state_4_3_63_32_sva_4
      & state_0_36_lpi_6) ^ (state_3_3_63_32_sva_4 & state_0_36_lpi_6);
  assign xor_cse_2030 = state_4_3_63_32_sva_11 & state_0_43_lpi_6;
  assign xor_cse_2029 = state_0_60_lpi_6 ^ xor_cse_1899 ^ xor_cse_1900 ^ xor_cse_2030;
  assign xor_cse_2032 = state_3_3_63_32_sva_11 & state_0_43_lpi_6;
  assign xor_cse_2033 = state_4_3_63_32_sva_5 ^ (state_4_3_63_32_sva_5 & state_0_37_lpi_6)
      ^ (state_3_3_63_32_sva_5 & state_0_37_lpi_6) ^ xor_cse_950;
  assign xor_cse_2036 = xor_cse_899 ^ state_4_3_63_32_sva_10 ^ (state_4_3_63_32_sva_10
      & state_0_42_lpi_6) ^ (state_3_3_63_32_sva_10 & state_0_42_lpi_6);
  assign xor_cse_2041 = state_4_3_63_32_sva_6 & state_0_38_lpi_6;
  assign xor_cse_2042 = state_3_3_63_32_sva_6 & state_0_38_lpi_6;
  assign xor_cse_2040 = xor_cse_2041 ^ xor_cse_2042 ^ state_4_3_63_32_sva_6;
  assign xor_cse_2045 = state_4_3_63_32_sva_9 & state_0_41_lpi_6;
  assign xor_cse_2046 = state_3_3_63_32_sva_9 & state_0_41_lpi_6;
  assign xor_cse_2044 = xor_cse_2045 ^ xor_cse_2046 ^ state_4_3_63_32_sva_9;
  assign xor_cse_2047 = xor_cse_867 ^ state_4_3_63_32_sva_7 ^ (state_4_3_63_32_sva_7
      & state_0_39_lpi_6) ^ (state_3_3_63_32_sva_7 & state_0_39_lpi_6);
  assign xor_cse_2054 = state_4_3_63_32_sva_8 & state_0_40_lpi_6;
  assign xor_cse_2055 = state_3_3_63_32_sva_8 & state_0_40_lpi_6;
  assign xor_cse_2053 = xor_cse_2054 ^ xor_cse_2055 ^ state_4_3_63_32_sva_8;
  assign xor_cse_2065 = xor_cse_2030 ^ xor_cse_2032 ^ state_4_3_63_32_sva_11;
  assign xor_cse_2069 = xor_cse_2022 ^ xor_cse_2024 ^ state_4_3_63_32_sva_12;
  assign xor_cse_2086 = xor_cse_107 ^ Encrypt_Top_sbox_1_and_596 ^ (state_3_39_lpi_3
      & state_1_1_63_32_lpi_4_7) ^ Encrypt_Top_sbox_1_and_1_cse_39_sva_1;
  assign xor_cse_2089 = state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_1_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_1_and_520 ^ (state_3_61_lpi_3 & state_1_1_63_32_lpi_4_29);
  assign xor_cse_2091 = AD_P6_AD_P6_xor_8_psp_sva_1 & state_3_0_lpi_3;
  assign xor_cse_2095 = ENC_P6_ENC_P6_xor_8_psp_sva_1 & state_3_0_lpi_3;
  assign xor_cse_2096 = xor_cse_164 ^ state_1_1_63_32_lpi_4_5 ^ Encrypt_Top_sbox_1_and_520
      ^ (state_3_61_lpi_3 & state_1_1_63_32_lpi_4_5);
  assign xor_cse_2098 = state_1_1_63_32_lpi_4_13 ^ xor_cse_107 ^ Encrypt_Top_sbox_1_and_596
      ^ (state_3_39_lpi_3 & state_1_1_63_32_lpi_4_13);
  assign xor_cse_2100 = xor_cse_196 ^ Encrypt_Top_sbox_1_and_628 ^ state_2_0_1_lpi_4
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[0]) ^ Encrypt_Top_sbox_3_and_1_cse_0_sva_1
      ^ (INIT_P12_INIT_P12_xor_8_psp_sva_1 & state_3_0_lpi_3);
  assign xor_cse_2104 = xor_cse_334 ^ (state_4_4_26_lpi_3 & state_0_26_lpi_6) ^ (state_3_26_lpi_3
      & state_0_26_lpi_6) ^ state_4_4_26_lpi_3;
  assign xor_cse_2106 = Encrypt_Top_sbox_2_and_648 ^ Encrypt_Top_sbox_2_and_650 ^
      state_4_4_16_lpi_3 ^ Encrypt_Top_sbox_2_and_756;
  assign state_3_16_sva_3_mx0w5 = xor_cse_2104 ^ xor_cse_242 ^ xor_cse_25 ^ xor_cse_2106
      ^ Encrypt_Top_sbox_2_and_758 ^ state_1_1_31_0_lpi_4_9;
  assign xor_cse_2109 = AD_P6_AD_P6_xor_7_psp_sva_1 & state_3_1_lpi_3;
  assign xor_cse_2108 = xor_cse_206 ^ Encrypt_Top_sbox_1_and_630 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ xor_cse_2109;
  assign xor_cse_2110 = state_2_1_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_1_sva_1;
  assign xor_cse_2112 = state_1_1_63_32_lpi_4_30 ^ Encrypt_Top_sbox_1_and_1_cse_62_sva_1
      ^ Encrypt_Top_sbox_1_and_518 ^ (state_3_62_lpi_3 & state_1_1_63_32_lpi_4_30);
  assign xor_cse_2113 = state_1_1_63_32_lpi_4_8 ^ Encrypt_Top_sbox_1_and_592 ^ (state_3_40_lpi_3
      & state_1_1_63_32_lpi_4_8) ^ Encrypt_Top_sbox_1_and_1_cse_40_sva_1;
  assign xor_cse_2111 = xor_cse_174 ^ xor_cse_120 ^ xor_cse_2112 ^ xor_cse_2113;
  assign xor_cse_2115 = ENC_P6_ENC_P6_xor_7_psp_sva_1 & state_3_1_lpi_3;
  assign xor_cse_2114 = xor_cse_206 ^ Encrypt_Top_sbox_1_and_630 ^ xor_cse_2115 ^
      state_2_1_1_lpi_6;
  assign xor_cse_2118 = xor_cse_120 ^ state_1_1_63_32_lpi_4_14 ^ Encrypt_Top_sbox_1_and_592
      ^ (state_3_40_lpi_3 & state_1_1_63_32_lpi_4_14);
  assign xor_cse_2120 = state_1_1_63_32_lpi_4_6 ^ xor_cse_174 ^ Encrypt_Top_sbox_1_and_518
      ^ (state_3_62_lpi_3 & state_1_1_63_32_lpi_4_6);
  assign xor_cse_2123 = state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[1])
      ^ Encrypt_Top_sbox_3_and_1_cse_1_sva_1 ^ (INIT_P12_INIT_P12_xor_7_psp_sva_1
      & state_3_1_lpi_3);
  assign xor_cse_2126 = xor_cse_38 ^ Encrypt_Top_sbox_2_and_750 ^ Encrypt_Top_sbox_2_and_748
      ^ Encrypt_Top_sbox_2_and_656;
  assign state_3_17_sva_3_mx0w5 = xor_cse_2126 ^ xor_cse_1317 ^ xor_cse_252 ^ Encrypt_Top_sbox_2_and_658
      ^ state_4_4_17_lpi_3 ^ state_1_1_63_32_lpi_4_0;
  assign xor_cse_2129 = xor_cse_217 ^ Encrypt_Top_sbox_1_and_632 ^ xor_cse_130 ^
      (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]);
  assign xor_cse_2131 = state_1_1_63_32_lpi_4_9 ^ Encrypt_Top_sbox_1_and_588 ^ (state_3_41_lpi_3
      & state_1_1_63_32_lpi_4_9) ^ Encrypt_Top_sbox_1_and_1_cse_41_sva_1;
  assign xor_cse_2132 = state_1_1_63_32_lpi_4_31 ^ Encrypt_Top_sbox_1_and_516 ^ (state_3_63_lpi_3
      & state_1_1_63_32_lpi_4_31) ^ Encrypt_Top_sbox_1_and_1_cse_63_sva_1;
  assign xor_cse_2134 = AD_P6_AD_P6_xor_6_psp_sva_1 & state_3_2_lpi_3;
  assign xor_cse_2137 = ENC_P6_ENC_P6_xor_6_psp_sva_1 & state_3_2_lpi_3;
  assign xor_cse_2138 = xor_cse_185 ^ state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_1_and_516
      ^ (state_3_63_lpi_3 & state_1_1_63_32_lpi_4_7);
  assign xor_cse_2142 = state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ Encrypt_Top_sbox_3_and_1_cse_2_sva_1 ^ (INIT_P12_INIT_P12_xor_6_psp_sva_1
      & state_3_2_lpi_3);
  assign xor_cse_2145 = state_3_41_lpi_3 & state_1_1_63_32_lpi_4_15;
  assign state_3_27_sva_3_mx0w5 = xor_cse_34 ^ xor_cse_1317 ^ xor_cse_80 ^ Encrypt_Top_sbox_2_and_724
      ^ Encrypt_Top_sbox_2_and_726 ^ state_1_1_63_32_lpi_4_11;
  assign xor_cse_2148 = xor_cse_196 ^ xor_cse_228 ^ xor_cse_8 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0])
      ^ Encrypt_Top_sbox_1_and_628 ^ Encrypt_Top_sbox_1_and_634 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]);
  assign xor_cse_2151 = state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_1_and_584 ^ (state_3_42_lpi_3
      & state_1_1_63_32_lpi_4_10) ^ Encrypt_Top_sbox_1_and_1_cse_42_sva_1;
  assign xor_cse_2153 = AD_P6_AD_P6_xor_5_psp_sva_1 & state_3_3_lpi_3;
  assign xor_cse_2157 = ENC_P6_ENC_P6_xor_5_psp_sva_1 & state_3_3_lpi_3;
  assign xor_cse_2159 = xor_cse_8 ^ state_1_1_63_32_lpi_4_16 ^ Encrypt_Top_sbox_1_and_584
      ^ (state_3_42_lpi_3 & state_1_1_63_32_lpi_4_16);
  assign xor_cse_2162 = state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ Encrypt_Top_sbox_3_and_1_cse_3_sva_1 ^ (INIT_P12_INIT_P12_xor_5_psp_sva_1
      & state_3_3_lpi_3);
  assign state_3_9_sva_3_mx0w5 = xor_cse_2104 ^ xor_cse_285 ^ xor_cse_274 ^ Encrypt_Top_sbox_2_and_672
      ^ Encrypt_Top_sbox_2_and_674 ^ state_4_4_19_lpi_3;
  assign xor_cse_2167 = xor_cse_22 ^ Encrypt_Top_sbox_1_and_580 ^ (state_3_43_lpi_3
      & state_1_1_63_32_lpi_4_11) ^ Encrypt_Top_sbox_1_and_1_cse_43_sva_1;
  assign xor_cse_2168 = xor_cse_206 ^ xor_cse_238 ^ state_1_1_63_32_lpi_4_11 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ Encrypt_Top_sbox_1_and_630 ^ Encrypt_Top_sbox_1_and_636 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign xor_cse_2172 = AD_P6_AD_P6_xor_4_psp_sva_1 & state_3_4_lpi_3;
  assign xor_cse_2176 = ENC_P6_ENC_P6_xor_4_psp_sva_1 & state_3_4_lpi_3;
  assign xor_cse_2178 = xor_cse_22 ^ state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_1_and_580
      ^ (state_3_43_lpi_3 & state_1_1_63_32_lpi_4_17);
  assign xor_cse_2182 = state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4])
      ^ Encrypt_Top_sbox_3_and_1_cse_4_sva_1 ^ (INIT_P12_INIT_P12_xor_4_psp_sva_1
      & state_3_4_lpi_3);
  assign xor_cse_2184 = xor_cse_102 ^ state_4_4_3_lpi_3 ^ state_4_4_37_lpi_3;
  assign state_4_60_sva_2_mx0w5 = xor_cse_2184 ^ state_1_1_63_32_lpi_4_11 ^ xor_cse_499
      ^ state_4_4_60_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_37_sva_1 ^ state_3_37_lpi_3
      ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1;
  assign xor_cse_2187 = state_1_1_63_32_lpi_4_12 ^ xor_cse_35 ^ Encrypt_Top_sbox_1_and_576
      ^ (state_3_44_lpi_3 & state_1_1_63_32_lpi_4_12);
  assign xor_cse_2190 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2]) ^ Encrypt_Top_sbox_1_and_632
      ^ Encrypt_Top_sbox_1_and_638 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]);
  assign xor_cse_2192 = AD_P6_AD_P6_xor_3_psp_sva_1 & state_3_5_lpi_3;
  assign xor_cse_2196 = ENC_P6_ENC_P6_xor_3_psp_sva_1 & state_3_5_lpi_3;
  assign xor_cse_2197 = xor_cse_248 ^ Encrypt_Top_sbox_1_and_638 ^ state_2_5_1_lpi_4
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[5]) ^ Encrypt_Top_sbox_3_and_1_cse_5_sva_1
      ^ (INIT_P12_INIT_P12_xor_3_psp_sva_1 & state_3_5_lpi_3);
  assign xor_cse_2201 = state_3_44_lpi_3 & state_1_1_63_32_lpi_4_18;
  assign state_4_61_sva_2_mx0w5 = xor_cse_111 ^ xor_cse_515 ^ xor_cse_588 ^ state_4_4_61_lpi_3
      ^ state_4_4_4_lpi_3 ^ state_4_4_38_lpi_3;
  assign xor_cse_2204 = xor_cse_49 ^ Encrypt_Top_sbox_1_and_572 ^ (state_3_45_lpi_3
      & state_1_1_63_32_lpi_4_13) ^ Encrypt_Top_sbox_1_and_1_cse_45_sva_1;
  assign xor_cse_2205 = xor_cse_258 ^ xor_cse_228 ^ state_1_1_63_32_lpi_4_13 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6])
      ^ Encrypt_Top_sbox_1_and_640 ^ Encrypt_Top_sbox_1_and_634 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]);
  assign xor_cse_2209 = AD_P6_AD_P6_xor_2_psp_sva_1 & state_3_6_lpi_3;
  assign xor_cse_2213 = ENC_P6_ENC_P6_xor_2_psp_sva_1 & state_3_6_lpi_3;
  assign xor_cse_2215 = state_1_1_63_32_lpi_4_19 ^ xor_cse_49 ^ Encrypt_Top_sbox_1_and_572
      ^ (state_3_45_lpi_3 & state_1_1_63_32_lpi_4_19);
  assign xor_cse_2219 = state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6])
      ^ Encrypt_Top_sbox_3_and_1_cse_6_sva_1 ^ (INIT_P12_INIT_P12_xor_2_psp_sva_1
      & state_3_6_lpi_3);
  assign xor_cse_2221 = xor_cse_124 ^ state_4_4_5_lpi_3 ^ state_4_4_39_lpi_3;
  assign state_4_62_sva_2_mx0w5 = xor_cse_2221 ^ state_1_1_63_32_lpi_4_13 ^ xor_cse_521
      ^ state_4_4_62_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_39_sva_1 ^ state_3_39_lpi_3
      ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1;
  assign xor_cse_2224 = xor_cse_63 ^ Encrypt_Top_sbox_1_and_568 ^ (state_3_46_lpi_3
      & state_1_1_63_32_lpi_4_14) ^ Encrypt_Top_sbox_1_and_1_cse_46_sva_1;
  assign xor_cse_2227 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]) ^ Encrypt_Top_sbox_1_and_642
      ^ Encrypt_Top_sbox_1_and_636 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign xor_cse_2229 = AD_P6_AD_P6_xor_1_psp_sva_1 & state_3_7_lpi_3;
  assign xor_cse_2230 = xor_cse_268 ^ (ENC_P6_ENC_P6_xor_1_psp_sva_1 & state_3_7_lpi_3)
      ^ state_2_7_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_7_sva_1;
  assign xor_cse_2234 = xor_cse_268 ^ Encrypt_Top_sbox_1_and_642 ^ state_2_7_1_lpi_4
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[7]) ^ Encrypt_Top_sbox_3_and_1_cse_7_sva_1
      ^ (INIT_P12_INIT_P12_xor_1_psp_sva_1 & state_3_7_lpi_3);
  assign xor_cse_2237 = state_1_1_63_32_lpi_4_2 ^ xor_cse_63 ^ Encrypt_Top_sbox_1_and_568
      ^ (state_3_46_lpi_3 & state_1_1_63_32_lpi_4_2);
  assign xor_cse_2241 = state_4_4_63_lpi_3 ^ state_4_4_6_lpi_3 ^ state_4_4_40_lpi_3;
  assign state_4_63_sva_2_mx0w5 = xor_cse_136 ^ xor_cse_527 ^ xor_cse_635 ^ xor_cse_2241;
  assign xor_cse_2242 = xor_cse_10 ^ Encrypt_Top_sbox_1_and_556 ^ (state_3_49_lpi_3
      & state_1_1_63_32_lpi_4_17) ^ Encrypt_Top_sbox_1_and_1_cse_49_sva_1;
  assign xor_cse_2243 = xor_cse_268 ^ Encrypt_Top_sbox_1_and_642 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7])
      ^ xor_cse_2229;
  assign xor_cse_2245 = state_4_4_10_lpi_3 ^ (state_2_10_1_lpi_4 & state_3_10_lpi_3)
      ^ (state_3_10_lpi_3 & state_1_1_31_0_lpi_4_10) ^ Encrypt_Top_sbox_1_and_1_cse_10_sva_1;
  assign xor_cse_2249 = state_1_1_63_32_lpi_4_22 ^ xor_cse_10 ^ Encrypt_Top_sbox_1_and_556
      ^ (state_3_49_lpi_3 & state_1_1_63_32_lpi_4_22);
  assign xor_cse_2252 = xor_cse_52 ^ Encrypt_Top_sbox_2_and_740 ^ Encrypt_Top_sbox_2_and_742
      ^ Encrypt_Top_sbox_2_and_664;
  assign state_3_18_sva_3_mx0w5 = xor_cse_1324 ^ xor_cse_2252 ^ xor_cse_263 ^ Encrypt_Top_sbox_2_and_666
      ^ state_4_4_18_lpi_3 ^ state_1_1_63_32_lpi_4_1;
  assign xor_cse_2255 = state_1_1_31_0_lpi_4_8 ^ Encrypt_Top_sbox_1_and_534 ^ (state_3_8_lpi_3
      & state_1_1_31_0_lpi_4_8) ^ Encrypt_Top_sbox_1_and_1_cse_8_sva_1;
  assign xor_cse_2256 = xor_cse_24 ^ Encrypt_Top_sbox_1_and_552 ^ (state_3_50_lpi_3
      & state_1_1_63_32_lpi_4_18) ^ Encrypt_Top_sbox_1_and_1_cse_50_sva_1;
  assign xor_cse_2258 = state_4_4_11_lpi_3 ^ (state_2_11_1_lpi_4 & state_3_11_lpi_3)
      ^ (state_3_11_lpi_3 & state_1_1_31_0_lpi_4_11) ^ Encrypt_Top_sbox_1_and_1_cse_11_sva_1;
  assign xor_cse_2259 = xor_cse_24 ^ state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_1_and_552
      ^ (state_3_50_lpi_3 & state_1_1_63_32_lpi_4_23);
  assign xor_cse_2262 = state_3_8_lpi_3 & state_1_1_63_32_lpi_4_8;
  assign xor_cse_2261 = Encrypt_Top_sbox_1_and_534 ^ xor_cse_2262 ^ Encrypt_Top_sbox_3_and_1_cse_8_sva_1
      ^ state_1_1_63_32_lpi_4_8;
  assign xor_cse_2264 = xor_cse_66 ^ Encrypt_Top_sbox_2_and_732 ^ Encrypt_Top_sbox_2_and_734
      ^ Encrypt_Top_sbox_2_and_672;
  assign xor_cse_2265 = xor_cse_274 ^ Encrypt_Top_sbox_2_and_674 ^ state_4_4_19_lpi_3
      ^ Encrypt_Top_sbox_2_and_752;
  assign state_3_19_sva_3_mx0w4 = xor_cse_2264 ^ xor_cse_2265 ^ xor_cse_369 ^ Encrypt_Top_sbox_2_and_754
      ^ state_4_4_29_lpi_3 ^ state_1_1_63_32_lpi_4_10;
  assign xor_cse_2268 = state_1_1_31_0_lpi_4_9 ^ Encrypt_Top_sbox_1_and_538 ^ (state_3_9_lpi_3
      & state_1_1_31_0_lpi_4_9) ^ Encrypt_Top_sbox_1_and_1_cse_9_sva_1;
  assign xor_cse_2269 = xor_cse_37 ^ Encrypt_Top_sbox_1_and_548 ^ (state_3_51_lpi_3
      & state_1_1_63_32_lpi_4_19) ^ Encrypt_Top_sbox_1_and_1_cse_51_sva_1;
  assign xor_cse_2271 = state_4_4_12_lpi_3 ^ (state_2_12_1_lpi_4 & state_3_12_lpi_3)
      ^ (state_3_12_lpi_3 & state_1_1_31_0_lpi_4_12) ^ Encrypt_Top_sbox_1_and_1_cse_12_sva_1;
  assign xor_cse_2272 = xor_cse_37 ^ state_1_1_63_32_lpi_4_24 ^ Encrypt_Top_sbox_1_and_548
      ^ (state_3_51_lpi_3 & state_1_1_63_32_lpi_4_24);
  assign xor_cse_2274 = xor_cse_286 ^ Encrypt_Top_sbox_1_and_538 ^ (state_3_9_lpi_3
      & state_1_1_63_32_lpi_4_9) ^ Encrypt_Top_sbox_3_and_1_cse_9_sva_1;
  assign xor_cse_2278 = state_4_4_19_lpi_3 ^ Encrypt_Top_sbox_2_and_672 ^ Encrypt_Top_sbox_2_and_674
      ^ Encrypt_Top_sbox_2_and_616;
  assign xor_cse_2279 = xor_cse_274 ^ Encrypt_Top_sbox_2_and_618 ^ state_4_4_12_lpi_3
      ^ xor_cse_204;
  assign state_3_2_sva_3_mx0w4 = xor_cse_217 ^ xor_cse_218 ^ xor_cse_2278 ^ xor_cse_2279;
  assign xor_cse_2280 = state_4_4_13_lpi_3 ^ (state_2_13_1_lpi_4 & state_3_13_lpi_3)
      ^ (state_3_13_lpi_3 & state_1_1_31_0_lpi_4_13) ^ Encrypt_Top_sbox_1_and_1_cse_13_sva_1;
  assign xor_cse_2281 = state_1_1_63_32_lpi_4_20 ^ xor_cse_51 ^ Encrypt_Top_sbox_1_and_544
      ^ (state_3_52_lpi_3 & state_1_1_63_32_lpi_4_20);
  assign xor_cse_2283 = xor_cse_51 ^ Encrypt_Top_sbox_1_and_544 ^ (state_3_52_lpi_3
      & state_1_1_63_32_lpi_4_25) ^ Encrypt_Top_sbox_3_and_1_cse_52_sva_1;
  assign xor_cse_2286 = xor_cse_80 ^ Encrypt_Top_sbox_2_and_724 ^ Encrypt_Top_sbox_2_and_726
      ^ Encrypt_Top_sbox_2_and_680;
  assign state_3_20_sva_3_mx0w4 = xor_cse_1341 ^ xor_cse_2286 ^ xor_cse_282 ^ Encrypt_Top_sbox_2_and_682
      ^ state_4_4_20_lpi_3 ^ state_1_1_63_32_lpi_4_11;
  assign xor_cse_2289 = xor_cse_221 ^ Encrypt_Top_sbox_1_and_1_cse_14_sva_1 ^ state_4_4_14_lpi_3
      ^ (state_2_14_1_lpi_4 & state_3_14_lpi_3);
  assign xor_cse_2290 = state_1_1_63_32_lpi_4_21 ^ xor_cse_65 ^ Encrypt_Top_sbox_1_and_540
      ^ (state_3_53_lpi_3 & state_1_1_63_32_lpi_4_21);
  assign xor_cse_2293 = xor_cse_65 ^ Encrypt_Top_sbox_1_and_540 ^ (state_3_53_lpi_3
      & state_1_1_63_32_lpi_4_26) ^ Encrypt_Top_sbox_3_and_1_cse_53_sva_1;
  assign xor_cse_2297 = state_1_1_63_32_lpi_4_12 ^ xor_cse_92 ^ Encrypt_Top_sbox_2_and_718
      ^ Encrypt_Top_sbox_2_and_716;
  assign state_3_21_sva_3_mx0w4 = xor_cse_2297 ^ xor_cse_1351 ^ xor_cse_1325;
  assign xor_cse_2298 = xor_cse_231 ^ Encrypt_Top_sbox_1_and_1_cse_15_sva_1 ^ state_4_4_15_lpi_3
      ^ (state_2_15_1_lpi_4 & state_3_15_lpi_3);
  assign xor_cse_2299 = xor_cse_79 ^ state_1_1_63_32_lpi_4_22 ^ Encrypt_Top_sbox_1_and_536
      ^ (state_3_54_lpi_3 & state_1_1_63_32_lpi_4_22);
  assign xor_cse_2302 = state_1_1_63_32_lpi_4_27 ^ xor_cse_79 ^ Encrypt_Top_sbox_1_and_536
      ^ (state_3_54_lpi_3 & state_1_1_63_32_lpi_4_27);
  assign state_3_22_sva_3_mx0w4 = xor_cse_1332 ^ xor_cse_1358 ^ xor_cse_107 ^ Encrypt_Top_sbox_2_and_708
      ^ Encrypt_Top_sbox_2_and_710 ^ state_1_1_63_32_lpi_4_13;
  assign xor_cse_2308 = xor_cse_242 ^ Encrypt_Top_sbox_1_and_1_cse_16_sva_1 ^ state_4_4_16_lpi_3
      ^ (state_2_16_1_lpi_4 & state_3_16_lpi_3);
  assign xor_cse_2309 = xor_cse_91 ^ Encrypt_Top_sbox_1_and_532 ^ (state_3_55_lpi_3
      & state_1_1_63_32_lpi_4_23) ^ Encrypt_Top_sbox_1_and_1_cse_55_sva_1;
  assign xor_cse_2313 = state_3_55_lpi_3 & state_1_1_63_32_lpi_4_28;
  assign xor_cse_2315 = xor_cse_25 ^ Encrypt_Top_sbox_2_and_758 ^ Encrypt_Top_sbox_2_and_756
      ^ Encrypt_Top_sbox_2_and_704;
  assign xor_cse_2316 = xor_cse_308 ^ Encrypt_Top_sbox_2_and_706 ^ state_4_4_23_lpi_3
      ^ Encrypt_Top_sbox_2_and_700;
  assign state_3_23_sva_3_mx0w4 = xor_cse_2315 ^ xor_cse_2316 ^ xor_cse_120 ^ state_1_1_31_0_lpi_4_9
      ^ Encrypt_Top_sbox_2_and_702 ^ state_1_1_63_32_lpi_4_14;
  assign xor_cse_2319 = xor_cse_106 ^ Encrypt_Top_sbox_1_and_530 ^ (state_3_56_lpi_3
      & state_1_1_63_32_lpi_4_24) ^ Encrypt_Top_sbox_1_and_1_cse_56_sva_1;
  assign xor_cse_2321 = Encrypt_Top_sbox_1_and_1_cse_17_sva_1 ^ state_4_4_17_lpi_3
      ^ (state_2_17_1_lpi_4 & state_3_17_lpi_3) ^ (state_3_17_lpi_3 & state_1_1_31_0_lpi_4_17);
  assign xor_cse_2323 = xor_cse_106 ^ Encrypt_Top_sbox_1_and_530 ^ (state_3_56_lpi_3
      & state_1_1_63_32_lpi_4_29) ^ Encrypt_Top_sbox_3_and_1_cse_56_sva_1;
  assign xor_cse_2327 = xor_cse_130 ^ Encrypt_Top_sbox_2_and_694 ^ Encrypt_Top_sbox_2_and_692
      ^ state_1_1_63_32_lpi_4_15;
  assign state_3_24_sva_3_mx0w4 = xor_cse_1350 ^ xor_cse_2327 ^ xor_cse_38 ^ Encrypt_Top_sbox_2_and_748
      ^ Encrypt_Top_sbox_2_and_750 ^ state_1_1_63_32_lpi_4_0;
  assign xor_cse_2331 = Encrypt_Top_sbox_1_and_1_cse_18_sva_1 ^ state_4_4_18_lpi_3
      ^ (state_2_18_1_lpi_4 & state_3_18_lpi_3) ^ (state_3_18_lpi_3 & state_1_1_31_0_lpi_4_18);
  assign xor_cse_2330 = xor_cse_263 ^ xor_cse_2331 ^ Encrypt_Top_sbox_1_and_654 ^
      Encrypt_Top_sbox_1_and_528;
  assign xor_cse_2333 = Encrypt_Top_sbox_1_and_728 ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1
      ^ state_1_1_63_32_lpi_4_25;
  assign xor_cse_2336 = state_3_57_lpi_3 & state_1_1_63_32_lpi_4_3;
  assign state_3_25_sva_3_mx0w4 = xor_cse_1357 ^ xor_cse_8 ^ xor_cse_52 ^ Encrypt_Top_sbox_2_and_740
      ^ Encrypt_Top_sbox_2_and_742 ^ state_1_1_63_32_lpi_4_1 ^ Encrypt_Top_sbox_2_and_684
      ^ Encrypt_Top_sbox_2_and_686 ^ state_1_1_63_32_lpi_4_16;
  assign xor_cse_2340 = xor_cse_132 ^ Encrypt_Top_sbox_1_and_526 ^ (state_3_58_lpi_3
      & state_1_1_63_32_lpi_4_26) ^ Encrypt_Top_sbox_1_and_1_cse_58_sva_1;
  assign xor_cse_2342 = Encrypt_Top_sbox_1_and_1_cse_19_sva_1 ^ state_4_4_19_lpi_3
      ^ (state_2_19_1_lpi_4 & state_3_19_lpi_3) ^ (state_3_19_lpi_3 & state_1_1_31_0_lpi_4_19);
  assign xor_cse_2344 = state_1_1_63_32_lpi_4_30 ^ xor_cse_132 ^ Encrypt_Top_sbox_1_and_526
      ^ (state_3_58_lpi_3 & state_1_1_63_32_lpi_4_30);
  assign state_3_26_sva_3_mx0w4 = xor_cse_2104 ^ xor_cse_22 ^ xor_cse_66 ^ Encrypt_Top_sbox_2_and_732
      ^ Encrypt_Top_sbox_2_and_734 ^ state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_2_and_676
      ^ Encrypt_Top_sbox_2_and_678 ^ state_1_1_63_32_lpi_4_17;
  assign xor_cse_2351 = xor_cse_282 ^ Encrypt_Top_sbox_1_and_1_cse_20_sva_1 ^ state_4_4_20_lpi_3
      ^ (state_2_20_1_lpi_4 & state_3_20_lpi_3);
  assign xor_cse_2352 = xor_cse_142 ^ Encrypt_Top_sbox_1_and_524 ^ (state_3_59_lpi_3
      & state_1_1_63_32_lpi_4_27) ^ Encrypt_Top_sbox_1_and_1_cse_59_sva_1;
  assign xor_cse_2356 = state_3_59_lpi_3 & state_1_1_63_32_lpi_4_31;
  assign state_3_28_sva_3_mx0w4 = xor_cse_2297 ^ xor_cse_1324 ^ xor_cse_49 ^ Encrypt_Top_sbox_2_and_660
      ^ Encrypt_Top_sbox_2_and_662 ^ state_1_1_63_32_lpi_4_19;
  assign xor_cse_2360 = xor_cse_290 ^ Encrypt_Top_sbox_1_and_1_cse_21_sva_1 ^ state_4_4_21_lpi_3
      ^ (state_2_21_1_lpi_4 & state_3_21_lpi_3);
  assign xor_cse_2361 = xor_cse_154 ^ Encrypt_Top_sbox_1_and_522 ^ Encrypt_Top_sbox_1_and_666
      ^ xor_cse_263;
  assign xor_cse_2366 = state_3_60_lpi_3 & state_1_1_63_32_lpi_4_4;
  assign xor_cse_2367 = xor_cse_107 ^ Encrypt_Top_sbox_2_and_710 ^ Encrypt_Top_sbox_2_and_708
      ^ Encrypt_Top_sbox_2_and_752;
  assign xor_cse_2370 = Encrypt_Top_sbox_2_and_654 ^ state_1_1_63_32_lpi_4_2;
  assign state_3_29_sva_3_mx0w4 = xor_cse_2367 ^ xor_cse_63 ^ xor_cse_369 ^ Encrypt_Top_sbox_2_and_754
      ^ state_4_4_29_lpi_3 ^ state_1_1_63_32_lpi_4_13 ^ Encrypt_Top_sbox_2_and_652
      ^ xor_cse_2370;
  assign xor_cse_2372 = state_4_4_22_lpi_3 ^ (state_2_22_1_lpi_4 & state_3_22_lpi_3)
      ^ (state_3_22_lpi_3 & state_1_1_31_0_lpi_4_22) ^ Encrypt_Top_sbox_1_and_1_cse_22_sva_1;
  assign xor_cse_2371 = xor_cse_299 ^ xor_cse_2372 ^ xor_cse_274 ^ xor_cse_2342;
  assign xor_cse_2373 = state_4_4_20_lpi_3 ^ Encrypt_Top_sbox_2_and_680 ^ Encrypt_Top_sbox_2_and_682
      ^ Encrypt_Top_sbox_2_and_624;
  assign xor_cse_2374 = xor_cse_282 ^ Encrypt_Top_sbox_2_and_626 ^ state_4_4_13_lpi_3
      ^ xor_cse_211;
  assign state_3_3_sva_3_mx0w4 = xor_cse_228 ^ xor_cse_229 ^ xor_cse_2373 ^ xor_cse_2374;
  assign xor_cse_2375 = state_4_4_23_lpi_3 ^ (state_2_23_1_lpi_4 & state_3_23_lpi_3)
      ^ (state_3_23_lpi_3 & state_1_1_31_0_lpi_4_23) ^ Encrypt_Top_sbox_1_and_1_cse_23_sva_1;
  assign xor_cse_2379 = xor_cse_120 ^ Encrypt_Top_sbox_2_and_700 ^ Encrypt_Top_sbox_2_and_702
      ^ Encrypt_Top_sbox_2_and_644;
  assign state_3_30_sva_3_mx0w4 = xor_cse_1341 ^ xor_cse_2379 ^ xor_cse_77 ^ state_1_1_63_32_lpi_4_14
      ^ Encrypt_Top_sbox_2_and_646 ^ state_1_1_63_32_lpi_4_20;
  assign xor_cse_2383 = state_4_4_24_lpi_3 ^ (state_2_24_1_lpi_4 & state_3_24_lpi_3)
      ^ (state_3_24_lpi_3 & state_1_1_31_0_lpi_4_24) ^ Encrypt_Top_sbox_1_and_1_cse_24_sva_1;
  assign xor_cse_2387 = Encrypt_Top_sbox_2_and_636 ^ Encrypt_Top_sbox_2_and_638 ^
      state_1_1_63_32_lpi_4_21;
  assign state_3_31_sva_3_mx0w4 = xor_cse_2327 ^ xor_cse_1351 ^ xor_cse_94 ^ xor_cse_2387;
  assign xor_cse_2388 = xor_cse_196 ^ Encrypt_Top_sbox_1_and_628 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0])
      ^ xor_cse_325;
  assign xor_cse_2390 = Encrypt_Top_sbox_1_and_1_cse_25_sva_1 ^ state_4_4_25_lpi_3
      ^ (state_2_25_1_lpi_4 & state_3_25_lpi_3) ^ (state_3_25_lpi_3 & state_1_1_31_0_lpi_4_25);
  assign xor_cse_2389 = xor_cse_299 ^ xor_cse_2372 ^ xor_cse_2390;
  assign xor_cse_2393 = state_4_4_21_lpi_3 ^ Encrypt_Top_sbox_2_and_688 ^ Encrypt_Top_sbox_2_and_690
      ^ Encrypt_Top_sbox_2_and_632;
  assign state_3_4_sva_3_mx0w5 = xor_cse_238 ^ xor_cse_221 ^ xor_cse_290 ^ xor_cse_239
      ^ xor_cse_2393 ^ Encrypt_Top_sbox_2_and_634 ^ state_4_4_14_lpi_3;
  assign xor_cse_2396 = state_4_4_26_lpi_3 ^ (state_2_26_1_lpi_4 & state_3_26_lpi_3)
      ^ (state_3_26_lpi_3 & state_1_1_31_0_lpi_4_26) ^ Encrypt_Top_sbox_1_and_1_cse_26_sva_1;
  assign xor_cse_2395 = xor_cse_308 ^ xor_cse_2375 ^ xor_cse_334 ^ xor_cse_2396;
  assign xor_cse_2397 = state_4_4_15_lpi_3 ^ Encrypt_Top_sbox_2_and_640 ^ Encrypt_Top_sbox_2_and_642
      ^ Encrypt_Top_sbox_2_and_696;
  assign xor_cse_2398 = xor_cse_231 ^ Encrypt_Top_sbox_2_and_698 ^ state_4_4_22_lpi_3
      ^ xor_cse_299;
  assign state_3_5_sva_3_mx0w5 = xor_cse_248 ^ xor_cse_249 ^ xor_cse_2397 ^ xor_cse_2398;
  assign xor_cse_2400 = state_4_4_27_lpi_3 ^ (state_2_27_1_lpi_4 & state_3_27_lpi_3)
      ^ (state_3_27_lpi_3 & state_1_1_31_0_lpi_4_27) ^ Encrypt_Top_sbox_1_and_1_cse_27_sva_1;
  assign xor_cse_2399 = xor_cse_343 ^ xor_cse_2400 ^ Encrypt_Top_sbox_1_and_632 ^
      xor_cse_217;
  assign xor_cse_2405 = state_4_4_16_lpi_3 ^ Encrypt_Top_sbox_2_and_648 ^ Encrypt_Top_sbox_2_and_650
      ^ Encrypt_Top_sbox_2_and_704;
  assign xor_cse_2406 = xor_cse_308 ^ Encrypt_Top_sbox_2_and_706 ^ state_4_4_23_lpi_3
      ^ xor_cse_242;
  assign state_3_6_sva_3_mx0w5 = xor_cse_258 ^ xor_cse_260 ^ xor_cse_2405 ^ xor_cse_2406;
  assign xor_cse_2408 = state_4_4_28_lpi_3 ^ (state_2_28_1_lpi_4 & state_3_28_lpi_3)
      ^ (state_3_28_lpi_3 & state_1_1_31_0_lpi_4_28) ^ Encrypt_Top_sbox_1_and_1_cse_28_sva_1;
  assign xor_cse_2407 = xor_cse_357 ^ xor_cse_2408 ^ Encrypt_Top_sbox_1_and_634 ^
      xor_cse_228;
  assign xor_cse_2413 = xor_cse_252 ^ Encrypt_Top_sbox_2_and_658 ^ state_4_4_17_lpi_3
      ^ Encrypt_Top_sbox_2_and_656;
  assign state_3_7_sva_3_mx0w5 = xor_cse_268 ^ xor_cse_270 ^ xor_cse_1350 ^ xor_cse_2413;
  assign xor_cse_2414 = xor_cse_238 ^ Encrypt_Top_sbox_1_and_636 ^ xor_cse_334 ^
      xor_cse_369;
  assign xor_cse_2416 = state_4_4_29_lpi_3 ^ (state_2_29_1_lpi_4 & state_3_29_lpi_3)
      ^ (state_3_29_lpi_3 & state_1_1_31_0_lpi_4_29) ^ Encrypt_Top_sbox_1_and_1_cse_29_sva_1;
  assign xor_cse_2421 = Encrypt_Top_sbox_2_and_664 ^ Encrypt_Top_sbox_2_and_666 ^
      state_4_4_18_lpi_3;
  assign state_3_8_sva_3_mx0w5 = xor_cse_1357 ^ xor_cse_277 ^ xor_cse_263 ^ xor_cse_2421;
  assign xor_cse_2422 = state_4_4_30_lpi_3 ^ (state_2_30_1_lpi_4 & state_3_30_lpi_3)
      ^ (state_3_30_lpi_3 & state_1_1_31_0_lpi_4_30) ^ Encrypt_Top_sbox_1_and_1_cse_30_sva_1;
  assign xor_cse_2423 = state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5])
      ^ Encrypt_Top_sbox_1_and_1_cse_5_sva_1 ^ xor_cse_2192;
  assign xor_cse_2426 = state_4_4_58_lpi_3 ^ state_4_4_1_lpi_3 ^ state_4_4_35_lpi_3;
  assign state_4_58_sva_2_mx0w5 = xor_cse_70 ^ xor_cse_480 ^ xor_cse_458 ^ xor_cse_2426;
  assign xor_cse_2427 = xor_cse_258 ^ Encrypt_Top_sbox_1_and_640 ^ xor_cse_357 ^
      xor_cse_394;
  assign xor_cse_2429 = state_4_4_31_lpi_3 ^ (state_2_31_1_lpi_4 & state_3_31_lpi_3)
      ^ (state_3_31_lpi_3 & state_1_1_31_0_lpi_4_31) ^ Encrypt_Top_sbox_1_and_1_cse_31_sva_1;
  assign state_4_59_sva_2_mx0w5 = xor_cse_84 ^ xor_cse_492 ^ state_4_4_59_lpi_3 ^
      state_4_4_2_lpi_3 ^ Encrypt_Top_sbox_3_and_cse_36_sva_1 ^ state_4_4_36_lpi_3
      ^ state_3_36_lpi_3 ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1 ^ state_1_1_63_32_lpi_4_10;
  assign xor_cse_2435 = state_1_1_63_32_lpi_4_15 ^ Encrypt_Top_sbox_1_and_564 ^ (state_3_47_lpi_3
      & state_1_1_63_32_lpi_4_15) ^ Encrypt_Top_sbox_1_and_1_cse_47_sva_1;
  assign xor_cse_2436 = xor_cse_248 ^ Encrypt_Top_sbox_1_and_638 ^ xor_cse_278 ^
      xor_cse_77;
  assign xor_cse_2439 = state_1_1_31_0_lpi_4_8 ^ xor_cse_11 ^ Encrypt_Top_sbox_1_and_624
      ^ (state_3_32_lpi_3 & state_1_1_31_0_lpi_4_8);
  assign xor_cse_2442 = xor_cse_258 ^ Encrypt_Top_sbox_1_and_640 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6])
      ^ Encrypt_Top_sbox_1_and_560;
  assign xor_cse_2443 = state_1_1_63_32_lpi_4_16 ^ (state_3_48_lpi_3 & state_1_1_63_32_lpi_4_16)
      ^ Encrypt_Top_sbox_1_and_1_cse_48_sva_1 ^ xor_cse_94;
  assign xor_cse_2448 = state_1_1_31_0_lpi_4_9 ^ xor_cse_25 ^ (state_3_33_lpi_3 &
      state_1_1_31_0_lpi_4_9) ^ Encrypt_Top_sbox_3_and_1_cse_33_sva_1;
  assign xor_cse_2452 = xor_cse_11 ^ Encrypt_Top_sbox_1_and_624 ^ (state_3_32_lpi_3
      & state_1_1_63_32_lpi_4_0) ^ Encrypt_Top_sbox_1_and_1_cse_32_sva_1;
  assign xor_cse_2457 = xor_cse_38 ^ Encrypt_Top_sbox_1_and_616 ^ (state_3_34_lpi_3
      & state_1_1_63_32_lpi_4_0) ^ Encrypt_Top_sbox_3_and_1_cse_34_sva_1;
  assign xor_cse_2461 = xor_cse_25 ^ state_1_1_63_32_lpi_4_1 ^ Encrypt_Top_sbox_1_and_694
      ^ Encrypt_Top_sbox_1_and_620;
  assign xor_cse_2463 = xor_cse_52 ^ Encrypt_Top_sbox_1_and_612 ^ (state_3_35_lpi_3
      & state_1_1_63_32_lpi_4_1) ^ Encrypt_Top_sbox_3_and_1_cse_35_sva_1;
  assign xor_cse_2468 = xor_cse_189 ^ xor_cse_2258 ^ Encrypt_Top_sbox_1_and_608 ^
      Encrypt_Top_sbox_1_and_620;
  assign xor_cse_2469 = state_1_1_63_32_lpi_4_10 ^ xor_cse_66 ^ (state_3_36_lpi_3
      & state_1_1_63_32_lpi_4_10) ^ Encrypt_Top_sbox_3_and_1_cse_36_sva_1;
  assign xor_cse_2472 = xor_cse_80 ^ Encrypt_Top_sbox_1_and_604 ^ (state_3_37_lpi_3
      & state_1_1_63_32_lpi_4_11) ^ Encrypt_Top_sbox_3_and_1_cse_37_sva_1;
  assign xor_cse_2476 = xor_cse_274 ^ xor_cse_2342 ^ xor_cse_130;
  assign xor_cse_2477 = xor_cse_92 ^ Encrypt_Top_sbox_1_and_600 ^ (state_3_38_lpi_3
      & state_1_1_63_32_lpi_4_12) ^ Encrypt_Top_sbox_3_and_1_cse_38_sva_1;
  assign xor_cse_2488 = Encrypt_Top_sbox_1_and_588 ^ xor_cse_2145 ^ Encrypt_Top_sbox_3_and_1_cse_41_sva_1
      ^ state_1_1_63_32_lpi_4_15;
  assign xor_cse_2505 = state_1_1_63_32_lpi_4_2 ^ xor_cse_38 ^ Encrypt_Top_sbox_1_and_616
      ^ (state_3_34_lpi_3 & state_1_1_63_32_lpi_4_2);
  assign xor_cse_2510 = state_1_1_63_32_lpi_4_20 ^ xor_cse_77 ^ Encrypt_Top_sbox_1_and_564
      ^ (state_3_47_lpi_3 & state_1_1_63_32_lpi_4_20);
  assign xor_cse_2516 = state_1_1_63_32_lpi_4_21 ^ xor_cse_94 ^ Encrypt_Top_sbox_1_and_560
      ^ (state_3_48_lpi_3 & state_1_1_63_32_lpi_4_21);
  assign xor_cse_2543 = xor_cse_119 ^ Encrypt_Top_sbox_1_and_528 ^ state_1_1_63_32_lpi_4_3
      ^ Encrypt_Top_sbox_1_and_522;
  assign xor_cse_2544 = xor_cse_52 ^ Encrypt_Top_sbox_1_and_612 ^ (state_3_35_lpi_3
      & state_1_1_63_32_lpi_4_3) ^ Encrypt_Top_sbox_1_and_1_cse_35_sva_1;
  assign xor_cse_2545 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1
      ^ Encrypt_Top_sbox_1_and_734 ^ xor_cse_154;
  assign xor_cse_2549 = state_1_1_63_32_lpi_4_4 ^ xor_cse_66 ^ (state_3_36_lpi_3
      & state_1_1_63_32_lpi_4_4) ^ Encrypt_Top_sbox_1_and_1_cse_36_sva_1;
  assign xor_cse_2559 = state_1_1_63_32_lpi_4_5 ^ xor_cse_80 ^ Encrypt_Top_sbox_1_and_604
      ^ (state_3_37_lpi_3 & state_1_1_63_32_lpi_4_5);
  assign xor_cse_2565 = state_1_1_63_32_lpi_4_6 ^ xor_cse_92 ^ Encrypt_Top_sbox_1_and_600
      ^ (state_3_38_lpi_3 & state_1_1_63_32_lpi_4_6);
  assign xor_cse_2598 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]) ^ Encrypt_Top_sbox_2_and_520
      ^ Encrypt_Top_sbox_2_and_522 ^ state_2_0_1_lpi_4;
  assign xor_cse_2602 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]) ^ Encrypt_Top_sbox_2_and_528
      ^ Encrypt_Top_sbox_2_and_530 ^ state_2_1_1_lpi_4;
  assign xor_cse_2604 = xor_cse_206 ^ state_2_1_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ Encrypt_Top_sbox_2_and_528;
  assign xor_cse_2608 = xor_cse_217 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2])
      ^ Encrypt_Top_sbox_2_and_536 ^ Encrypt_Top_sbox_2_and_538;
  assign xor_cse_2610 = xor_cse_228 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3])
      ^ Encrypt_Top_sbox_2_and_544 ^ Encrypt_Top_sbox_2_and_546;
  assign xor_cse_2612 = xor_cse_238 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4])
      ^ Encrypt_Top_sbox_2_and_552 ^ Encrypt_Top_sbox_2_and_554;
  assign xor_cse_2618 = xor_cse_248 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5])
      ^ Encrypt_Top_sbox_2_and_560 ^ Encrypt_Top_sbox_2_and_562;
  assign xor_cse_2620 = xor_cse_258 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6])
      ^ Encrypt_Top_sbox_2_and_568 ^ Encrypt_Top_sbox_2_and_570;
  assign xor_cse_2625 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]) ^ Encrypt_Top_sbox_2_and_576
      ^ Encrypt_Top_sbox_2_and_578 ^ state_2_7_1_lpi_6;
  assign xor_cse_2626 = state_1_1_63_32_lpi_4_9 ^ state_4_4_41_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_41_sva_1
      ^ state_3_41_lpi_3;
  assign state_4_0_sva_3 = xor_cse_148 ^ xor_cse_56 ^ xor_cse_643 ^ state_4_4_0_lpi_3
      ^ state_4_4_7_lpi_3 ^ state_1_1_63_32_lpi_4_15;
  assign xor_cse_2629 = state_1_1_63_32_lpi_4_10 ^ state_4_4_42_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_42_sva_1
      ^ state_3_42_lpi_3;
  assign state_4_1_sva_3 = xor_cse_70 ^ xor_cse_587 ^ xor_cse_651 ^ state_4_4_1_lpi_3
      ^ state_4_4_8_lpi_3 ^ state_4_4_42_lpi_3;
  assign xor_cse_2641 = state_1_1_63_32_lpi_4_0 ^ Encrypt_Top_sbox_2_and_764 ^ xor_cse_11
      ^ Encrypt_Top_sbox_2_and_766;
  assign xor_cse_2688 = state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_2_and_668 ^ Encrypt_Top_sbox_2_and_670
      ^ xor_cse_35;
  assign xor_cse_2707 = xor_cse_94 ^ Encrypt_Top_sbox_2_and_636 ^ Encrypt_Top_sbox_2_and_638
      ^ state_1_1_63_32_lpi_4_16;
  assign xor_cse_2771 = xor_cse_132 ^ Encrypt_Top_sbox_2_and_558 ^ state_1_1_63_32_lpi_4_26
      ^ Encrypt_Top_sbox_2_and_556;
  assign xor_cse_2791 = xor_cse_174 ^ Encrypt_Top_sbox_2_and_526 ^ state_1_1_63_32_lpi_4_30;
  assign xor_cse_2799 = xor_cse_185 ^ Encrypt_Top_sbox_2_and_518 ^ state_1_1_63_32_lpi_4_31;
  assign xor_cse_2808 = xor_cse_196 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0])
      ^ state_2_0_1_lpi_6 ^ Encrypt_Top_sbox_2_and_520;
  assign xor_cse_2814 = state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_2_and_628 ^ Encrypt_Top_sbox_2_and_630
      ^ Encrypt_Top_sbox_2_and_548;
  assign xor_cse_2822 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_2_and_542 ^ Encrypt_Top_sbox_2_and_540
      ^ Encrypt_Top_sbox_2_and_620;
  assign xor_cse_2827 = state_1_1_63_32_lpi_4_19 ^ xor_cse_37 ^ state_1_1_63_32_lpi_4_29
      ^ xor_cse_164;
  assign xor_cse_2830 = state_1_1_63_32_lpi_4_20 ^ Encrypt_Top_sbox_2_and_604 ^ Encrypt_Top_sbox_2_and_606
      ^ Encrypt_Top_sbox_2_and_524;
  assign xor_cse_2836 = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6]) ^ Encrypt_Top_sbox_2_and_568
      ^ Encrypt_Top_sbox_2_and_570 ^ Encrypt_Top_sbox_2_and_596;
  assign xor_cse_2848 = state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_2_and_580 ^ Encrypt_Top_sbox_2_and_582
      ^ Encrypt_Top_sbox_2_and_584;
  assign xor_cse_2855 = state_1_1_31_0_lpi_4_9 ^ Encrypt_Top_sbox_2_and_592 ^ Encrypt_Top_sbox_2_and_594
      ^ Encrypt_Top_sbox_2_and_572;
  assign xor_cse_2868 = xor_cse_278 ^ Encrypt_Top_sbox_2_and_586 ^ state_1_1_31_0_lpi_4_8
      ^ Encrypt_Top_sbox_2_and_584;
  assign xor_cse_2887 = state_1_1_31_0_lpi_4_10 ^ Encrypt_Top_sbox_2_and_2_cse_17_sva_1
      ^ state_4_4_51_lpi_3;
  assign state_4_10_sva_3 = xor_cse_479 ^ xor_cse_717 ^ xor_cse_569 ^ xor_cse_2887;
  assign xor_cse_2889 = Encrypt_Top_sbox_2_and_2_cse_11_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1
      ^ state_4_4_52_lpi_3;
  assign state_4_11_sva_3 = xor_cse_594 ^ xor_cse_491 ^ xor_cse_726 ^ xor_cse_2889;
  assign xor_cse_2891 = Encrypt_Top_sbox_2_and_2_cse_12_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1
      ^ state_4_4_53_lpi_3;
  assign state_4_12_sva_3 = xor_cse_603 ^ xor_cse_498 ^ xor_cse_734 ^ xor_cse_2891;
  assign xor_cse_2893 = Encrypt_Top_sbox_2_and_2_cse_13_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1
      ^ state_4_4_54_lpi_3;
  assign state_4_13_sva_3 = xor_cse_609 ^ xor_cse_514 ^ xor_cse_740 ^ xor_cse_2893;
  assign xor_cse_2895 = Encrypt_Top_sbox_2_and_2_cse_14_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1
      ^ state_4_4_55_lpi_3;
  assign state_4_14_sva_3 = xor_cse_618 ^ xor_cse_520 ^ xor_cse_746 ^ xor_cse_2895;
  assign xor_cse_2897 = Encrypt_Top_sbox_2_and_2_cse_15_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_22_sva_1
      ^ state_4_4_56_lpi_3;
  assign state_4_15_sva_3 = xor_cse_673 ^ xor_cse_752 ^ xor_cse_528 ^ xor_cse_2897;
  assign xor_cse_2903 = state_1_1_63_32_lpi_4_27 ^ Encrypt_Top_sbox_1_and_cse_59_sva_1
      ^ state_4_4_59_lpi_3 ^ state_3_59_lpi_3;
  assign xor_cse_2906 = state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_2_and_2_cse_60_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_60_sva_1 ^ state_4_4_60_lpi_3;
  assign xor_cse_2909 = state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_2_and_2_cse_61_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_61_sva_1 ^ state_4_4_61_lpi_3;
  assign xor_cse_2912 = state_4_4_62_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_62_sva_1
      ^ state_3_62_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_62_sva_1;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      data_out_rsci_idat_0 <= 1'b0;
      data_out_rsci_idat_1 <= 1'b0;
      data_out_rsci_idat_2 <= 1'b0;
      data_out_rsci_idat_3 <= 1'b0;
      data_out_rsci_idat_4 <= 1'b0;
      data_out_rsci_idat_5 <= 1'b0;
      data_out_rsci_idat_6 <= 1'b0;
      data_out_rsci_idat_7 <= 1'b0;
      data_out_rsci_idat_8 <= 1'b0;
      data_out_rsci_idat_9 <= 1'b0;
      data_out_rsci_idat_10 <= 1'b0;
      data_out_rsci_idat_11 <= 1'b0;
      data_out_rsci_idat_12 <= 1'b0;
      data_out_rsci_idat_13 <= 1'b0;
      data_out_rsci_idat_14 <= 1'b0;
      data_out_rsci_idat_15 <= 1'b0;
      data_out_rsci_idat_16 <= 1'b0;
      data_out_rsci_idat_17 <= 1'b0;
      data_out_rsci_idat_18 <= 1'b0;
      data_out_rsci_idat_19 <= 1'b0;
      data_out_rsci_idat_20 <= 1'b0;
      data_out_rsci_idat_21 <= 1'b0;
      data_out_rsci_idat_22 <= 1'b0;
      data_out_rsci_idat_23 <= 1'b0;
      data_out_rsci_idat_24 <= 1'b0;
      data_out_rsci_idat_25 <= 1'b0;
      data_out_rsci_idat_26 <= 1'b0;
      data_out_rsci_idat_27 <= 1'b0;
      data_out_rsci_idat_28 <= 1'b0;
      data_out_rsci_idat_29 <= 1'b0;
      data_out_rsci_idat_30 <= 1'b0;
      data_out_rsci_idat_31 <= 1'b0;
    end
    else if ( rst ) begin
      data_out_rsci_idat_0 <= 1'b0;
      data_out_rsci_idat_1 <= 1'b0;
      data_out_rsci_idat_2 <= 1'b0;
      data_out_rsci_idat_3 <= 1'b0;
      data_out_rsci_idat_4 <= 1'b0;
      data_out_rsci_idat_5 <= 1'b0;
      data_out_rsci_idat_6 <= 1'b0;
      data_out_rsci_idat_7 <= 1'b0;
      data_out_rsci_idat_8 <= 1'b0;
      data_out_rsci_idat_9 <= 1'b0;
      data_out_rsci_idat_10 <= 1'b0;
      data_out_rsci_idat_11 <= 1'b0;
      data_out_rsci_idat_12 <= 1'b0;
      data_out_rsci_idat_13 <= 1'b0;
      data_out_rsci_idat_14 <= 1'b0;
      data_out_rsci_idat_15 <= 1'b0;
      data_out_rsci_idat_16 <= 1'b0;
      data_out_rsci_idat_17 <= 1'b0;
      data_out_rsci_idat_18 <= 1'b0;
      data_out_rsci_idat_19 <= 1'b0;
      data_out_rsci_idat_20 <= 1'b0;
      data_out_rsci_idat_21 <= 1'b0;
      data_out_rsci_idat_22 <= 1'b0;
      data_out_rsci_idat_23 <= 1'b0;
      data_out_rsci_idat_24 <= 1'b0;
      data_out_rsci_idat_25 <= 1'b0;
      data_out_rsci_idat_26 <= 1'b0;
      data_out_rsci_idat_27 <= 1'b0;
      data_out_rsci_idat_28 <= 1'b0;
      data_out_rsci_idat_29 <= 1'b0;
      data_out_rsci_idat_30 <= 1'b0;
      data_out_rsci_idat_31 <= 1'b0;
    end
    else if ( and_4636_cse ) begin
      data_out_rsci_idat_0 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_2_itm_mx0w0, state_0_0_sva_2_mx0w1,
          ciphertext_32_sva_mx0w2, PLEN_xor_62_nl, xor_403_nl, xor_262_nl, data_out_rsci_idat_0_mx0w6,
          data_out_rsci_idat_0_mx0w7, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse
          , (fsm_output[12]) , and_94_cse , (fsm_output[15]) , (fsm_output[16]) ,
          (fsm_output[17])});
      data_out_rsci_idat_1 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_4_itm_mx0w0, state_0_1_sva_2_mx0w1,
          ciphertext_33_sva_mx0w2, PLEN_xor_60_nl, xor_418_nl, xor_260_nl, data_out_rsci_idat_1_mx0w6,
          data_out_rsci_idat_1_mx0w7, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse
          , (fsm_output[12]) , and_94_cse , (fsm_output[15]) , (fsm_output[16]) ,
          (fsm_output[17])});
      data_out_rsci_idat_2 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_6_itm_mx0w0, state_0_2_sva_2_mx0w1,
          ciphertext_34_sva_mx0w2, PLEN_xor_58_nl, xor_432_nl, xor_258_nl, data_out_rsci_idat_2_mx0w6,
          xor_321_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_3 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_8_itm_mx0w0, state_0_3_sva_2_mx0w1,
          ciphertext_35_sva_mx0w2, PLEN_xor_56_nl, xor_447_nl, xor_256_nl, data_out_rsci_idat_3_mx0w6,
          xor_319_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_4 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_10_itm_mx0w0, state_0_4_sva_2_mx0w1,
          ciphertext_36_sva_mx0w2, PLEN_xor_54_nl, xor_462_nl, xor_254_nl, data_out_rsci_idat_4_mx0w6,
          xor_317_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_5 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_12_itm_mx0w0, state_0_5_sva_2_mx0w1,
          ciphertext_37_sva_mx0w2, PLEN_xor_52_nl, xor_477_nl, xor_252_nl, data_out_rsci_idat_5_mx0w6,
          xor_315_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_6 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_14_itm_mx0w0, state_0_6_sva_2_mx0w1,
          ciphertext_38_sva_mx0w2, PLEN_xor_50_nl, xor_492_nl, xor_250_nl, data_out_rsci_idat_6_mx0w6,
          xor_313_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_7 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_16_itm_mx0w0, state_0_7_sva_2_mx0w1,
          ciphertext_39_sva_mx0w2, PLEN_xor_48_nl, xor_506_nl, xor_248_nl, data_out_rsci_idat_7_mx0w6,
          xor_311_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_8 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_18_itm_mx0w0, state_0_8_sva_2_mx0w1,
          ciphertext_40_sva_mx0w2, PLEN_xor_46_nl, xor_520_nl, xor_246_nl, data_out_rsci_idat_8_mx0w6,
          data_out_rsci_idat_8_mx0w7, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse
          , (fsm_output[12]) , and_94_cse , (fsm_output[15]) , (fsm_output[16]) ,
          (fsm_output[17])});
      data_out_rsci_idat_9 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_20_itm_mx0w0, state_0_9_sva_2_mx0w1,
          ciphertext_41_sva_mx0w2, PLEN_xor_44_nl, xor_533_nl, xor_244_nl, data_out_rsci_idat_9_mx0w6,
          data_out_rsci_idat_9_mx0w7, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse
          , (fsm_output[12]) , and_94_cse , (fsm_output[15]) , (fsm_output[16]) ,
          (fsm_output[17])});
      data_out_rsci_idat_10 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_22_itm_mx0w0, state_0_10_sva_2_mx0w1,
          ciphertext_42_sva_mx0w2, PLEN_xor_42_nl, xor_546_nl, xor_242_nl, data_out_rsci_idat_10_mx0w6,
          xor_305_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_11 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_24_itm_mx0w0, state_0_11_sva_2_mx0w1,
          ciphertext_43_sva_mx0w2, PLEN_xor_40_nl, xor_558_nl, xor_240_nl, data_out_rsci_idat_11_mx0w6,
          xor_303_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_12 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_26_itm_mx0w0, state_0_12_sva_2_mx0w1,
          ciphertext_44_sva_mx0w2, PLEN_xor_38_nl, xor_568_nl, xor_238_nl, data_out_rsci_idat_12_mx0w6,
          xor_301_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_13 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_28_itm_mx0w0, state_0_13_sva_2_mx0w1,
          ciphertext_45_sva_mx0w2, PLEN_xor_36_nl, xor_579_nl, xor_236_nl, data_out_rsci_idat_13_mx0w6,
          xor_299_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_14 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_30_itm_mx0w0, state_0_14_sva_2_mx0w1,
          ciphertext_46_sva_mx0w2, PLEN_xor_34_nl, xor_591_nl, xor_234_nl, data_out_rsci_idat_14_mx0w6,
          xor_297_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_15 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_32_itm_mx0w0, state_0_15_sva_2_mx0w1,
          ciphertext_47_sva_mx0w2, PLEN_xor_nl, xor_604_nl, xor_232_nl, data_out_rsci_idat_15_mx0w6,
          xor_295_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_16 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_34_itm_mx0w0, state_0_16_sva_2_mx0w1,
          ciphertext_48_sva_mx0w2, PLEN_xor_33_nl, xor_615_nl, xor_230_nl, data_out_rsci_idat_16_mx0w6,
          xor_293_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_17 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_36_itm_mx0w0, state_0_17_sva_2_mx0w1,
          ciphertext_49_sva_mx0w2, PLEN_xor_35_nl, xor_626_nl, xor_228_nl, data_out_rsci_idat_17_mx0w6,
          xor_291_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_18 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_38_itm_mx0w0, state_0_18_sva_2_mx0w1,
          ciphertext_50_sva_mx0w2, PLEN_xor_37_nl, xor_637_nl, xor_226_nl, data_out_rsci_idat_18_mx0w6,
          xor_289_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_19 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_40_itm_mx0w0, state_0_19_sva_2_mx0w1,
          ciphertext_51_sva_mx0w2, PLEN_xor_39_nl, xor_649_nl, xor_224_nl, data_out_rsci_idat_19_mx0w6,
          xor_287_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_20 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_42_itm_mx0w0, state_0_20_sva_2_mx0w1,
          ciphertext_52_sva_mx0w2, PLEN_xor_41_nl, xor_660_nl, xor_222_nl, data_out_rsci_idat_20_mx0w6,
          xor_285_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_21 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_44_itm_mx0w0, state_0_21_sva_2_mx0w1,
          ciphertext_53_sva_mx0w2, PLEN_xor_43_nl, xor_672_nl, xor_220_nl, data_out_rsci_idat_21_mx0w6,
          xor_283_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_22 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_46_itm_mx0w0, state_0_22_sva_2_mx0w1,
          ciphertext_54_sva_mx0w2, PLEN_xor_45_nl, xor_683_nl, xor_218_nl, data_out_rsci_idat_22_mx0w6,
          xor_281_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_23 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_48_itm_mx0w0, state_0_23_sva_2_mx0w1,
          ciphertext_55_sva_mx0w2, PLEN_xor_47_nl, xor_692_nl, xor_216_nl, data_out_rsci_idat_23_mx0w6,
          xor_279_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_24 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_50_itm_mx0w0, state_0_24_sva_2_mx0w1,
          ciphertext_56_sva_mx0w2, PLEN_xor_49_nl, xor_701_nl, xor_214_nl, data_out_rsci_idat_24_mx0w6,
          xor_277_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_25 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_52_itm_mx0w0, state_0_25_sva_2_mx0w1,
          ciphertext_57_sva_mx0w2, PLEN_xor_51_nl, xor_711_nl, xor_212_nl, data_out_rsci_idat_25_mx0w6,
          xor_275_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_26 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_54_itm_mx0w0, state_0_26_sva_2_mx0w1,
          ciphertext_58_sva_mx0w2, PLEN_xor_53_nl, xor_721_nl, xor_210_nl, xor_316_nl,
          xor_273_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_27 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_56_itm_mx0w0, state_0_27_sva_2_mx0w1,
          ciphertext_59_sva_mx0w2, PLEN_xor_55_nl, xor_731_nl, xor_208_nl, xor_318_nl,
          xor_271_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_28 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_58_itm_mx0w0, state_0_28_sva_2_mx0w1,
          ciphertext_60_sva_mx0w2, PLEN_xor_57_nl, xor_741_nl, xor_206_nl, xor_320_nl,
          xor_269_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_29 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_60_itm_mx0w0, state_0_29_sva_2_mx0w1,
          ciphertext_61_sva_mx0w2, PLEN_xor_59_nl, xor_751_nl, xor_204_nl, xor_322_nl,
          xor_267_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_30 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_62_itm_mx0w0, state_0_30_sva_2_mx0w1,
          ciphertext_62_sva_mx0w2, PLEN_xor_61_nl, xor_760_nl, xor_202_nl, xor_324_nl,
          xor_265_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
      data_out_rsci_idat_31 <= MUX1HOT_s_1_8_2(ADLEN_ADLEN_xor_64_itm_mx0w0, state_0_31_sva_2_mx0w1,
          ciphertext_63_sva_mx0w2, PLEN_xor_63_nl, xor_769_nl, xor_9_nl, xor_326_nl,
          xor_11_nl, {(fsm_output[6]) , (fsm_output[7]) , and_90_cse , (fsm_output[12])
          , and_94_cse , (fsm_output[15]) , (fsm_output[16]) , (fsm_output[17])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_4_3_63_32_sva_31 <= 1'b0;
      state_4_3_63_32_sva_30 <= 1'b0;
      state_4_3_63_32_sva_29 <= 1'b0;
      state_4_3_63_32_sva_28 <= 1'b0;
      state_4_3_63_32_sva_27 <= 1'b0;
      state_4_3_63_32_sva_26 <= 1'b0;
      state_4_3_63_32_sva_25 <= 1'b0;
      state_4_3_63_32_sva_24 <= 1'b0;
      state_4_3_63_32_sva_23 <= 1'b0;
      state_4_3_63_32_sva_22 <= 1'b0;
      state_4_3_63_32_sva_21 <= 1'b0;
      state_4_3_63_32_sva_20 <= 1'b0;
      state_4_3_63_32_sva_19 <= 1'b0;
      state_4_3_63_32_sva_18 <= 1'b0;
      state_4_3_63_32_sva_17 <= 1'b0;
      state_4_3_63_32_sva_16 <= 1'b0;
      state_4_3_63_32_sva_15 <= 1'b0;
      state_4_3_63_32_sva_14 <= 1'b0;
      state_4_3_63_32_sva_13 <= 1'b0;
      state_4_3_63_32_sva_12 <= 1'b0;
      state_4_3_63_32_sva_11 <= 1'b0;
      state_4_3_63_32_sva_10 <= 1'b0;
      state_4_3_63_32_sva_9 <= 1'b0;
      state_4_3_63_32_sva_8 <= 1'b0;
      state_4_3_63_32_sva_7 <= 1'b0;
      state_4_3_63_32_sva_6 <= 1'b0;
      state_4_3_63_32_sva_5 <= 1'b0;
      state_4_3_63_32_sva_4 <= 1'b0;
      state_4_3_63_32_sva_3 <= 1'b0;
      state_4_3_63_32_sva_2 <= 1'b0;
      state_4_3_63_32_sva_1 <= 1'b0;
      state_4_3_63_32_sva_0 <= 1'b0;
      state_3_3_63_32_sva_31 <= 1'b0;
      state_3_3_63_32_sva_30 <= 1'b0;
      state_3_3_63_32_sva_29 <= 1'b0;
      state_3_3_63_32_sva_28 <= 1'b0;
      state_3_3_63_32_sva_27 <= 1'b0;
      state_3_3_63_32_sva_26 <= 1'b0;
      state_3_3_63_32_sva_25 <= 1'b0;
      state_3_3_63_32_sva_24 <= 1'b0;
      state_3_3_63_32_sva_23 <= 1'b0;
      state_3_3_63_32_sva_22 <= 1'b0;
      state_3_3_63_32_sva_21 <= 1'b0;
      state_3_3_63_32_sva_20 <= 1'b0;
      state_3_3_63_32_sva_19 <= 1'b0;
      state_3_3_63_32_sva_18 <= 1'b0;
      state_3_3_63_32_sva_17 <= 1'b0;
      state_3_3_63_32_sva_16 <= 1'b0;
      state_3_3_63_32_sva_15 <= 1'b0;
      state_3_3_63_32_sva_14 <= 1'b0;
      state_3_3_63_32_sva_13 <= 1'b0;
      state_3_3_63_32_sva_12 <= 1'b0;
      state_3_3_63_32_sva_11 <= 1'b0;
      state_3_3_63_32_sva_10 <= 1'b0;
      state_3_3_63_32_sva_9 <= 1'b0;
      state_3_3_63_32_sva_8 <= 1'b0;
      state_3_3_63_32_sva_7 <= 1'b0;
      state_3_3_63_32_sva_6 <= 1'b0;
      state_3_3_63_32_sva_5 <= 1'b0;
      state_3_3_63_32_sva_4 <= 1'b0;
      state_3_3_63_32_sva_3 <= 1'b0;
      state_3_3_63_32_sva_2 <= 1'b0;
      state_3_3_63_32_sva_1 <= 1'b0;
      state_3_3_63_32_sva_0 <= 1'b0;
      state_4_3_31_0_sva_31 <= 1'b0;
      state_4_3_31_0_sva_30 <= 1'b0;
      state_4_3_31_0_sva_29 <= 1'b0;
      state_4_3_31_0_sva_28 <= 1'b0;
      state_4_3_31_0_sva_27 <= 1'b0;
      state_4_3_31_0_sva_26 <= 1'b0;
      state_4_3_31_0_sva_25 <= 1'b0;
      state_4_3_31_0_sva_24 <= 1'b0;
      state_4_3_31_0_sva_23 <= 1'b0;
      state_4_3_31_0_sva_22 <= 1'b0;
      state_4_3_31_0_sva_21 <= 1'b0;
      state_4_3_31_0_sva_20 <= 1'b0;
      state_4_3_31_0_sva_19 <= 1'b0;
      state_4_3_31_0_sva_18 <= 1'b0;
      state_4_3_31_0_sva_17 <= 1'b0;
      state_4_3_31_0_sva_16 <= 1'b0;
      state_4_3_31_0_sva_15 <= 1'b0;
      state_4_3_31_0_sva_14 <= 1'b0;
      state_4_3_31_0_sva_13 <= 1'b0;
      state_4_3_31_0_sva_12 <= 1'b0;
      state_4_3_31_0_sva_11 <= 1'b0;
      state_4_3_31_0_sva_10 <= 1'b0;
      state_4_3_31_0_sva_9 <= 1'b0;
      state_4_3_31_0_sva_8 <= 1'b0;
      state_4_3_31_0_sva_7 <= 1'b0;
      state_4_3_31_0_sva_6 <= 1'b0;
      state_4_3_31_0_sva_5 <= 1'b0;
      state_4_3_31_0_sva_4 <= 1'b0;
      state_4_3_31_0_sva_3 <= 1'b0;
      state_4_3_31_0_sva_2 <= 1'b0;
      state_4_3_31_0_sva_1 <= 1'b0;
      state_4_3_31_0_sva_0 <= 1'b0;
      state_3_3_31_0_sva_31 <= 1'b0;
      state_3_3_31_0_sva_30 <= 1'b0;
      state_3_3_31_0_sva_29 <= 1'b0;
      state_3_3_31_0_sva_28 <= 1'b0;
      state_3_3_31_0_sva_27 <= 1'b0;
      state_3_3_31_0_sva_26 <= 1'b0;
      state_3_3_31_0_sva_25 <= 1'b0;
      state_3_3_31_0_sva_24 <= 1'b0;
      state_3_3_31_0_sva_23 <= 1'b0;
      state_3_3_31_0_sva_22 <= 1'b0;
      state_3_3_31_0_sva_21 <= 1'b0;
      state_3_3_31_0_sva_20 <= 1'b0;
      state_3_3_31_0_sva_19 <= 1'b0;
      state_3_3_31_0_sva_18 <= 1'b0;
      state_3_3_31_0_sva_17 <= 1'b0;
      state_3_3_31_0_sva_16 <= 1'b0;
      state_3_3_31_0_sva_15 <= 1'b0;
      state_3_3_31_0_sva_14 <= 1'b0;
      state_3_3_31_0_sva_13 <= 1'b0;
      state_3_3_31_0_sva_12 <= 1'b0;
      state_3_3_31_0_sva_11 <= 1'b0;
      state_3_3_31_0_sva_10 <= 1'b0;
      state_3_3_31_0_sva_9 <= 1'b0;
      state_3_3_31_0_sva_8 <= 1'b0;
      state_3_3_31_0_sva_7 <= 1'b0;
      state_3_3_31_0_sva_6 <= 1'b0;
      state_3_3_31_0_sva_5 <= 1'b0;
      state_3_3_31_0_sva_4 <= 1'b0;
      state_3_3_31_0_sva_3 <= 1'b0;
      state_3_3_31_0_sva_2 <= 1'b0;
      state_3_3_31_0_sva_1 <= 1'b0;
      state_3_3_31_0_sva_0 <= 1'b0;
      reg_data_out_rsci_iswt0_cse <= 1'b0;
      reg_data_in_rsci_iswt0_cse <= 1'b0;
      AD_P6_j_2_0_sva <= 3'b000;
    end
    else if ( rst ) begin
      state_4_3_63_32_sva_31 <= 1'b0;
      state_4_3_63_32_sva_30 <= 1'b0;
      state_4_3_63_32_sva_29 <= 1'b0;
      state_4_3_63_32_sva_28 <= 1'b0;
      state_4_3_63_32_sva_27 <= 1'b0;
      state_4_3_63_32_sva_26 <= 1'b0;
      state_4_3_63_32_sva_25 <= 1'b0;
      state_4_3_63_32_sva_24 <= 1'b0;
      state_4_3_63_32_sva_23 <= 1'b0;
      state_4_3_63_32_sva_22 <= 1'b0;
      state_4_3_63_32_sva_21 <= 1'b0;
      state_4_3_63_32_sva_20 <= 1'b0;
      state_4_3_63_32_sva_19 <= 1'b0;
      state_4_3_63_32_sva_18 <= 1'b0;
      state_4_3_63_32_sva_17 <= 1'b0;
      state_4_3_63_32_sva_16 <= 1'b0;
      state_4_3_63_32_sva_15 <= 1'b0;
      state_4_3_63_32_sva_14 <= 1'b0;
      state_4_3_63_32_sva_13 <= 1'b0;
      state_4_3_63_32_sva_12 <= 1'b0;
      state_4_3_63_32_sva_11 <= 1'b0;
      state_4_3_63_32_sva_10 <= 1'b0;
      state_4_3_63_32_sva_9 <= 1'b0;
      state_4_3_63_32_sva_8 <= 1'b0;
      state_4_3_63_32_sva_7 <= 1'b0;
      state_4_3_63_32_sva_6 <= 1'b0;
      state_4_3_63_32_sva_5 <= 1'b0;
      state_4_3_63_32_sva_4 <= 1'b0;
      state_4_3_63_32_sva_3 <= 1'b0;
      state_4_3_63_32_sva_2 <= 1'b0;
      state_4_3_63_32_sva_1 <= 1'b0;
      state_4_3_63_32_sva_0 <= 1'b0;
      state_3_3_63_32_sva_31 <= 1'b0;
      state_3_3_63_32_sva_30 <= 1'b0;
      state_3_3_63_32_sva_29 <= 1'b0;
      state_3_3_63_32_sva_28 <= 1'b0;
      state_3_3_63_32_sva_27 <= 1'b0;
      state_3_3_63_32_sva_26 <= 1'b0;
      state_3_3_63_32_sva_25 <= 1'b0;
      state_3_3_63_32_sva_24 <= 1'b0;
      state_3_3_63_32_sva_23 <= 1'b0;
      state_3_3_63_32_sva_22 <= 1'b0;
      state_3_3_63_32_sva_21 <= 1'b0;
      state_3_3_63_32_sva_20 <= 1'b0;
      state_3_3_63_32_sva_19 <= 1'b0;
      state_3_3_63_32_sva_18 <= 1'b0;
      state_3_3_63_32_sva_17 <= 1'b0;
      state_3_3_63_32_sva_16 <= 1'b0;
      state_3_3_63_32_sva_15 <= 1'b0;
      state_3_3_63_32_sva_14 <= 1'b0;
      state_3_3_63_32_sva_13 <= 1'b0;
      state_3_3_63_32_sva_12 <= 1'b0;
      state_3_3_63_32_sva_11 <= 1'b0;
      state_3_3_63_32_sva_10 <= 1'b0;
      state_3_3_63_32_sva_9 <= 1'b0;
      state_3_3_63_32_sva_8 <= 1'b0;
      state_3_3_63_32_sva_7 <= 1'b0;
      state_3_3_63_32_sva_6 <= 1'b0;
      state_3_3_63_32_sva_5 <= 1'b0;
      state_3_3_63_32_sva_4 <= 1'b0;
      state_3_3_63_32_sva_3 <= 1'b0;
      state_3_3_63_32_sva_2 <= 1'b0;
      state_3_3_63_32_sva_1 <= 1'b0;
      state_3_3_63_32_sva_0 <= 1'b0;
      state_4_3_31_0_sva_31 <= 1'b0;
      state_4_3_31_0_sva_30 <= 1'b0;
      state_4_3_31_0_sva_29 <= 1'b0;
      state_4_3_31_0_sva_28 <= 1'b0;
      state_4_3_31_0_sva_27 <= 1'b0;
      state_4_3_31_0_sva_26 <= 1'b0;
      state_4_3_31_0_sva_25 <= 1'b0;
      state_4_3_31_0_sva_24 <= 1'b0;
      state_4_3_31_0_sva_23 <= 1'b0;
      state_4_3_31_0_sva_22 <= 1'b0;
      state_4_3_31_0_sva_21 <= 1'b0;
      state_4_3_31_0_sva_20 <= 1'b0;
      state_4_3_31_0_sva_19 <= 1'b0;
      state_4_3_31_0_sva_18 <= 1'b0;
      state_4_3_31_0_sva_17 <= 1'b0;
      state_4_3_31_0_sva_16 <= 1'b0;
      state_4_3_31_0_sva_15 <= 1'b0;
      state_4_3_31_0_sva_14 <= 1'b0;
      state_4_3_31_0_sva_13 <= 1'b0;
      state_4_3_31_0_sva_12 <= 1'b0;
      state_4_3_31_0_sva_11 <= 1'b0;
      state_4_3_31_0_sva_10 <= 1'b0;
      state_4_3_31_0_sva_9 <= 1'b0;
      state_4_3_31_0_sva_8 <= 1'b0;
      state_4_3_31_0_sva_7 <= 1'b0;
      state_4_3_31_0_sva_6 <= 1'b0;
      state_4_3_31_0_sva_5 <= 1'b0;
      state_4_3_31_0_sva_4 <= 1'b0;
      state_4_3_31_0_sva_3 <= 1'b0;
      state_4_3_31_0_sva_2 <= 1'b0;
      state_4_3_31_0_sva_1 <= 1'b0;
      state_4_3_31_0_sva_0 <= 1'b0;
      state_3_3_31_0_sva_31 <= 1'b0;
      state_3_3_31_0_sva_30 <= 1'b0;
      state_3_3_31_0_sva_29 <= 1'b0;
      state_3_3_31_0_sva_28 <= 1'b0;
      state_3_3_31_0_sva_27 <= 1'b0;
      state_3_3_31_0_sva_26 <= 1'b0;
      state_3_3_31_0_sva_25 <= 1'b0;
      state_3_3_31_0_sva_24 <= 1'b0;
      state_3_3_31_0_sva_23 <= 1'b0;
      state_3_3_31_0_sva_22 <= 1'b0;
      state_3_3_31_0_sva_21 <= 1'b0;
      state_3_3_31_0_sva_20 <= 1'b0;
      state_3_3_31_0_sva_19 <= 1'b0;
      state_3_3_31_0_sva_18 <= 1'b0;
      state_3_3_31_0_sva_17 <= 1'b0;
      state_3_3_31_0_sva_16 <= 1'b0;
      state_3_3_31_0_sva_15 <= 1'b0;
      state_3_3_31_0_sva_14 <= 1'b0;
      state_3_3_31_0_sva_13 <= 1'b0;
      state_3_3_31_0_sva_12 <= 1'b0;
      state_3_3_31_0_sva_11 <= 1'b0;
      state_3_3_31_0_sva_10 <= 1'b0;
      state_3_3_31_0_sva_9 <= 1'b0;
      state_3_3_31_0_sva_8 <= 1'b0;
      state_3_3_31_0_sva_7 <= 1'b0;
      state_3_3_31_0_sva_6 <= 1'b0;
      state_3_3_31_0_sva_5 <= 1'b0;
      state_3_3_31_0_sva_4 <= 1'b0;
      state_3_3_31_0_sva_3 <= 1'b0;
      state_3_3_31_0_sva_2 <= 1'b0;
      state_3_3_31_0_sva_1 <= 1'b0;
      state_3_3_31_0_sva_0 <= 1'b0;
      reg_data_out_rsci_iswt0_cse <= 1'b0;
      reg_data_in_rsci_iswt0_cse <= 1'b0;
      AD_P6_j_2_0_sva <= 3'b000;
    end
    else if ( run_wen ) begin
      state_4_3_63_32_sva_31 <= MUX_s_1_2_2((nonce3[31]), state_xor_338_nl, fsm_output[1]);
      state_4_3_63_32_sva_30 <= MUX_s_1_2_2((nonce3[30]), state_xor_340_nl, fsm_output[1]);
      state_4_3_63_32_sva_29 <= MUX_s_1_2_2((nonce3[29]), state_xor_342_nl, fsm_output[1]);
      state_4_3_63_32_sva_28 <= MUX_s_1_2_2((nonce3[28]), state_xor_344_nl, fsm_output[1]);
      state_4_3_63_32_sva_27 <= MUX_s_1_2_2((nonce3[27]), state_xor_346_nl, fsm_output[1]);
      state_4_3_63_32_sva_26 <= MUX_s_1_2_2((nonce3[26]), state_xor_348_nl, fsm_output[1]);
      state_4_3_63_32_sva_25 <= MUX_s_1_2_2((nonce3[25]), state_xor_350_nl, fsm_output[1]);
      state_4_3_63_32_sva_24 <= MUX_s_1_2_2((nonce3[24]), state_xor_352_nl, fsm_output[1]);
      state_4_3_63_32_sva_23 <= MUX_s_1_2_2((nonce3[23]), state_xor_354_nl, fsm_output[1]);
      state_4_3_63_32_sva_22 <= MUX_s_1_2_2((nonce3[22]), state_xor_356_nl, fsm_output[1]);
      state_4_3_63_32_sva_21 <= MUX_s_1_2_2((nonce3[21]), state_xor_358_nl, fsm_output[1]);
      state_4_3_63_32_sva_20 <= MUX_s_1_2_2((nonce3[20]), state_xor_360_nl, fsm_output[1]);
      state_4_3_63_32_sva_19 <= MUX_s_1_2_2((nonce3[19]), state_xor_362_nl, fsm_output[1]);
      state_4_3_63_32_sva_18 <= MUX_s_1_2_2((nonce3[18]), state_xor_364_nl, fsm_output[1]);
      state_4_3_63_32_sva_17 <= MUX_s_1_2_2((nonce3[17]), state_xor_366_nl, fsm_output[1]);
      state_4_3_63_32_sva_16 <= MUX_s_1_2_2((nonce3[16]), state_xor_368_nl, fsm_output[1]);
      state_4_3_63_32_sva_15 <= MUX_s_1_2_2((nonce3[15]), state_xor_370_nl, fsm_output[1]);
      state_4_3_63_32_sva_14 <= MUX_s_1_2_2((nonce3[14]), state_xor_372_nl, fsm_output[1]);
      state_4_3_63_32_sva_13 <= MUX_s_1_2_2((nonce3[13]), state_xor_374_nl, fsm_output[1]);
      state_4_3_63_32_sva_12 <= MUX_s_1_2_2((nonce3[12]), state_xor_376_nl, fsm_output[1]);
      state_4_3_63_32_sva_11 <= MUX_s_1_2_2((nonce3[11]), state_xor_378_nl, fsm_output[1]);
      state_4_3_63_32_sva_10 <= MUX_s_1_2_2((nonce3[10]), state_xor_380_nl, fsm_output[1]);
      state_4_3_63_32_sva_9 <= MUX_s_1_2_2((nonce3[9]), state_xor_382_nl, fsm_output[1]);
      state_4_3_63_32_sva_8 <= MUX_s_1_2_2((nonce3[8]), state_xor_384_nl, fsm_output[1]);
      state_4_3_63_32_sva_7 <= MUX_s_1_2_2((nonce3[7]), state_xor_386_nl, fsm_output[1]);
      state_4_3_63_32_sva_6 <= MUX_s_1_2_2((nonce3[6]), state_xor_388_nl, fsm_output[1]);
      state_4_3_63_32_sva_5 <= MUX_s_1_2_2((nonce3[5]), state_xor_390_nl, fsm_output[1]);
      state_4_3_63_32_sva_4 <= MUX_s_1_2_2((nonce3[4]), state_xor_392_nl, fsm_output[1]);
      state_4_3_63_32_sva_3 <= MUX_s_1_2_2((nonce3[3]), state_xor_394_nl, fsm_output[1]);
      state_4_3_63_32_sva_2 <= MUX_s_1_2_2((nonce3[2]), state_xor_396_nl, fsm_output[1]);
      state_4_3_63_32_sva_1 <= MUX_s_1_2_2((nonce3[1]), state_xor_398_nl, fsm_output[1]);
      state_4_3_63_32_sva_0 <= MUX_s_1_2_2((nonce3[0]), state_xor_400_nl, fsm_output[1]);
      state_3_3_63_32_sva_31 <= MUX_s_1_2_2((nonce1[31]), state_xor_402_nl, fsm_output[1]);
      state_3_3_63_32_sva_30 <= MUX_s_1_2_2((nonce1[30]), state_xor_404_nl, fsm_output[1]);
      state_3_3_63_32_sva_29 <= MUX_s_1_2_2((nonce1[29]), state_xor_406_nl, fsm_output[1]);
      state_3_3_63_32_sva_28 <= MUX_s_1_2_2((nonce1[28]), state_xor_408_nl, fsm_output[1]);
      state_3_3_63_32_sva_27 <= MUX_s_1_2_2((nonce1[27]), state_xor_410_nl, fsm_output[1]);
      state_3_3_63_32_sva_26 <= MUX_s_1_2_2((nonce1[26]), state_xor_412_nl, fsm_output[1]);
      state_3_3_63_32_sva_25 <= MUX_s_1_2_2((nonce1[25]), state_xor_414_nl, fsm_output[1]);
      state_3_3_63_32_sva_24 <= MUX_s_1_2_2((nonce1[24]), state_xor_416_nl, fsm_output[1]);
      state_3_3_63_32_sva_23 <= MUX_s_1_2_2((nonce1[23]), state_xor_418_nl, fsm_output[1]);
      state_3_3_63_32_sva_22 <= MUX_s_1_2_2((nonce1[22]), state_xor_420_nl, fsm_output[1]);
      state_3_3_63_32_sva_21 <= MUX_s_1_2_2((nonce1[21]), state_xor_422_nl, fsm_output[1]);
      state_3_3_63_32_sva_20 <= MUX_s_1_2_2((nonce1[20]), state_xor_424_nl, fsm_output[1]);
      state_3_3_63_32_sva_19 <= MUX_s_1_2_2((nonce1[19]), state_xor_426_nl, fsm_output[1]);
      state_3_3_63_32_sva_18 <= MUX_s_1_2_2((nonce1[18]), state_xor_428_nl, fsm_output[1]);
      state_3_3_63_32_sva_17 <= MUX_s_1_2_2((nonce1[17]), state_xor_430_nl, fsm_output[1]);
      state_3_3_63_32_sva_16 <= MUX_s_1_2_2((nonce1[16]), state_xor_432_nl, fsm_output[1]);
      state_3_3_63_32_sva_15 <= MUX_s_1_2_2((nonce1[15]), state_xor_434_nl, fsm_output[1]);
      state_3_3_63_32_sva_14 <= MUX_s_1_2_2((nonce1[14]), state_xor_436_nl, fsm_output[1]);
      state_3_3_63_32_sva_13 <= MUX_s_1_2_2((nonce1[13]), state_xor_438_nl, fsm_output[1]);
      state_3_3_63_32_sva_12 <= MUX_s_1_2_2((nonce1[12]), state_xor_440_nl, fsm_output[1]);
      state_3_3_63_32_sva_11 <= MUX_s_1_2_2((nonce1[11]), state_xor_442_nl, fsm_output[1]);
      state_3_3_63_32_sva_10 <= MUX_s_1_2_2((nonce1[10]), state_xor_444_nl, fsm_output[1]);
      state_3_3_63_32_sva_9 <= MUX_s_1_2_2((nonce1[9]), state_xor_446_nl, fsm_output[1]);
      state_3_3_63_32_sva_8 <= MUX_s_1_2_2((nonce1[8]), state_xor_448_nl, fsm_output[1]);
      state_3_3_63_32_sva_7 <= MUX_s_1_2_2((nonce1[7]), state_xor_450_nl, fsm_output[1]);
      state_3_3_63_32_sva_6 <= MUX_s_1_2_2((nonce1[6]), state_xor_452_nl, fsm_output[1]);
      state_3_3_63_32_sva_5 <= MUX_s_1_2_2((nonce1[5]), state_xor_454_nl, fsm_output[1]);
      state_3_3_63_32_sva_4 <= MUX_s_1_2_2((nonce1[4]), state_xor_456_nl, fsm_output[1]);
      state_3_3_63_32_sva_3 <= MUX_s_1_2_2((nonce1[3]), state_xor_458_nl, fsm_output[1]);
      state_3_3_63_32_sva_2 <= MUX_s_1_2_2((nonce1[2]), state_xor_460_nl, fsm_output[1]);
      state_3_3_63_32_sva_1 <= MUX_s_1_2_2((nonce1[1]), state_xor_462_nl, fsm_output[1]);
      state_3_3_63_32_sva_0 <= MUX_s_1_2_2((nonce1[0]), state_xor_464_nl, fsm_output[1]);
      state_4_3_31_0_sva_31 <= MUX_s_1_2_2((nonce4[31]), state_xor_401_nl, fsm_output[1]);
      state_4_3_31_0_sva_30 <= MUX_s_1_2_2((nonce4[30]), state_xor_399_nl, fsm_output[1]);
      state_4_3_31_0_sva_29 <= MUX_s_1_2_2((nonce4[29]), state_xor_397_nl, fsm_output[1]);
      state_4_3_31_0_sva_28 <= MUX_s_1_2_2((nonce4[28]), state_xor_395_nl, fsm_output[1]);
      state_4_3_31_0_sva_27 <= MUX_s_1_2_2((nonce4[27]), state_xor_393_nl, fsm_output[1]);
      state_4_3_31_0_sva_26 <= MUX_s_1_2_2((nonce4[26]), state_xor_391_nl, fsm_output[1]);
      state_4_3_31_0_sva_25 <= MUX_s_1_2_2((nonce4[25]), state_xor_389_nl, fsm_output[1]);
      state_4_3_31_0_sva_24 <= MUX_s_1_2_2((nonce4[24]), state_xor_387_nl, fsm_output[1]);
      state_4_3_31_0_sva_23 <= MUX_s_1_2_2((nonce4[23]), state_xor_385_nl, fsm_output[1]);
      state_4_3_31_0_sva_22 <= MUX_s_1_2_2((nonce4[22]), state_xor_383_nl, fsm_output[1]);
      state_4_3_31_0_sva_21 <= MUX_s_1_2_2((nonce4[21]), state_xor_381_nl, fsm_output[1]);
      state_4_3_31_0_sva_20 <= MUX_s_1_2_2((nonce4[20]), state_xor_379_nl, fsm_output[1]);
      state_4_3_31_0_sva_19 <= MUX_s_1_2_2((nonce4[19]), state_xor_377_nl, fsm_output[1]);
      state_4_3_31_0_sva_18 <= MUX_s_1_2_2((nonce4[18]), state_xor_375_nl, fsm_output[1]);
      state_4_3_31_0_sva_17 <= MUX_s_1_2_2((nonce4[17]), state_xor_373_nl, fsm_output[1]);
      state_4_3_31_0_sva_16 <= MUX_s_1_2_2((nonce4[16]), state_xor_371_nl, fsm_output[1]);
      state_4_3_31_0_sva_15 <= MUX_s_1_2_2((nonce4[15]), state_xor_369_nl, fsm_output[1]);
      state_4_3_31_0_sva_14 <= MUX_s_1_2_2((nonce4[14]), state_xor_367_nl, fsm_output[1]);
      state_4_3_31_0_sva_13 <= MUX_s_1_2_2((nonce4[13]), state_xor_365_nl, fsm_output[1]);
      state_4_3_31_0_sva_12 <= MUX_s_1_2_2((nonce4[12]), state_xor_363_nl, fsm_output[1]);
      state_4_3_31_0_sva_11 <= MUX_s_1_2_2((nonce4[11]), state_xor_361_nl, fsm_output[1]);
      state_4_3_31_0_sva_10 <= MUX_s_1_2_2((nonce4[10]), state_xor_359_nl, fsm_output[1]);
      state_4_3_31_0_sva_9 <= MUX_s_1_2_2((nonce4[9]), state_xor_357_nl, fsm_output[1]);
      state_4_3_31_0_sva_8 <= MUX_s_1_2_2((nonce4[8]), state_xor_355_nl, fsm_output[1]);
      state_4_3_31_0_sva_7 <= MUX_s_1_2_2((nonce4[7]), state_xor_353_nl, fsm_output[1]);
      state_4_3_31_0_sva_6 <= MUX_s_1_2_2((nonce4[6]), state_xor_351_nl, fsm_output[1]);
      state_4_3_31_0_sva_5 <= MUX_s_1_2_2((nonce4[5]), state_xor_349_nl, fsm_output[1]);
      state_4_3_31_0_sva_4 <= MUX_s_1_2_2((nonce4[4]), state_xor_347_nl, fsm_output[1]);
      state_4_3_31_0_sva_3 <= MUX_s_1_2_2((nonce4[3]), state_xor_345_nl, fsm_output[1]);
      state_4_3_31_0_sva_2 <= MUX_s_1_2_2((nonce4[2]), state_xor_343_nl, fsm_output[1]);
      state_4_3_31_0_sva_1 <= MUX_s_1_2_2((nonce4[1]), state_xor_341_nl, fsm_output[1]);
      state_4_3_31_0_sva_0 <= MUX_s_1_2_2((nonce4[0]), state_xor_339_nl, fsm_output[1]);
      state_3_3_31_0_sva_31 <= MUX_s_1_2_2((nonce2[31]), state_xor_465_nl, fsm_output[1]);
      state_3_3_31_0_sva_30 <= MUX_s_1_2_2((nonce2[30]), state_xor_463_nl, fsm_output[1]);
      state_3_3_31_0_sva_29 <= MUX_s_1_2_2((nonce2[29]), state_xor_461_nl, fsm_output[1]);
      state_3_3_31_0_sva_28 <= MUX_s_1_2_2((nonce2[28]), state_xor_459_nl, fsm_output[1]);
      state_3_3_31_0_sva_27 <= MUX_s_1_2_2((nonce2[27]), state_xor_457_nl, fsm_output[1]);
      state_3_3_31_0_sva_26 <= MUX_s_1_2_2((nonce2[26]), state_xor_455_nl, fsm_output[1]);
      state_3_3_31_0_sva_25 <= MUX_s_1_2_2((nonce2[25]), state_xor_453_nl, fsm_output[1]);
      state_3_3_31_0_sva_24 <= MUX_s_1_2_2((nonce2[24]), state_xor_451_nl, fsm_output[1]);
      state_3_3_31_0_sva_23 <= MUX_s_1_2_2((nonce2[23]), state_xor_449_nl, fsm_output[1]);
      state_3_3_31_0_sva_22 <= MUX_s_1_2_2((nonce2[22]), state_xor_447_nl, fsm_output[1]);
      state_3_3_31_0_sva_21 <= MUX_s_1_2_2((nonce2[21]), state_xor_445_nl, fsm_output[1]);
      state_3_3_31_0_sva_20 <= MUX_s_1_2_2((nonce2[20]), state_xor_443_nl, fsm_output[1]);
      state_3_3_31_0_sva_19 <= MUX_s_1_2_2((nonce2[19]), state_xor_441_nl, fsm_output[1]);
      state_3_3_31_0_sva_18 <= MUX_s_1_2_2((nonce2[18]), state_xor_439_nl, fsm_output[1]);
      state_3_3_31_0_sva_17 <= MUX_s_1_2_2((nonce2[17]), state_xor_437_nl, fsm_output[1]);
      state_3_3_31_0_sva_16 <= MUX_s_1_2_2((nonce2[16]), state_xor_435_nl, fsm_output[1]);
      state_3_3_31_0_sva_15 <= MUX_s_1_2_2((nonce2[15]), state_xor_433_nl, fsm_output[1]);
      state_3_3_31_0_sva_14 <= MUX_s_1_2_2((nonce2[14]), state_xor_431_nl, fsm_output[1]);
      state_3_3_31_0_sva_13 <= MUX_s_1_2_2((nonce2[13]), state_xor_429_nl, fsm_output[1]);
      state_3_3_31_0_sva_12 <= MUX_s_1_2_2((nonce2[12]), state_xor_427_nl, fsm_output[1]);
      state_3_3_31_0_sva_11 <= MUX_s_1_2_2((nonce2[11]), state_xor_425_nl, fsm_output[1]);
      state_3_3_31_0_sva_10 <= MUX_s_1_2_2((nonce2[10]), state_xor_423_nl, fsm_output[1]);
      state_3_3_31_0_sva_9 <= MUX_s_1_2_2((nonce2[9]), state_xor_421_nl, fsm_output[1]);
      state_3_3_31_0_sva_8 <= MUX_s_1_2_2((nonce2[8]), state_xor_419_nl, fsm_output[1]);
      state_3_3_31_0_sva_7 <= MUX_s_1_2_2((nonce2[7]), state_xor_417_nl, fsm_output[1]);
      state_3_3_31_0_sva_6 <= MUX_s_1_2_2((nonce2[6]), state_xor_415_nl, fsm_output[1]);
      state_3_3_31_0_sva_5 <= MUX_s_1_2_2((nonce2[5]), state_xor_413_nl, fsm_output[1]);
      state_3_3_31_0_sva_4 <= MUX_s_1_2_2((nonce2[4]), state_xor_411_nl, fsm_output[1]);
      state_3_3_31_0_sva_3 <= MUX_s_1_2_2((nonce2[3]), state_xor_409_nl, fsm_output[1]);
      state_3_3_31_0_sva_2 <= MUX_s_1_2_2((nonce2[2]), state_xor_407_nl, fsm_output[1]);
      state_3_3_31_0_sva_1 <= MUX_s_1_2_2((nonce2[1]), state_xor_405_nl, fsm_output[1]);
      state_3_3_31_0_sva_0 <= MUX_s_1_2_2((nonce2[0]), state_xor_403_nl, fsm_output[1]);
      reg_data_out_rsci_iswt0_cse <= or_2210_cse;
      reg_data_in_rsci_iswt0_cse <= and_738_cse | (fsm_output[2]) | (fsm_output[9])
          | (fsm_output[8]) | (fsm_output[6]) | (fsm_output[5]) | and_740_cse;
      AD_P6_j_2_0_sva <= MUX_v_3_2_2(3'b000, AD_P6_j_2_0_sva_2, and_24_cse);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_0_lpi_6 <= 1'b0;
      state_0_1_lpi_6 <= 1'b0;
      state_0_2_lpi_6 <= 1'b0;
      state_0_3_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_0_lpi_6 <= 1'b0;
      state_0_1_lpi_6 <= 1'b0;
      state_0_2_lpi_6 <= 1'b0;
      state_0_3_lpi_6 <= 1'b0;
    end
    else if ( state_and_cse ) begin
      state_0_0_lpi_6 <= mux1h_nl & (~ (fsm_output[0]));
      state_0_1_lpi_6 <= mux1h_1_nl & (~ (fsm_output[0]));
      state_0_2_lpi_6 <= mux1h_2_nl & (~ (fsm_output[0]));
      state_0_3_lpi_6 <= mux1h_3_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_4_lpi_6 <= 1'b0;
      state_0_5_lpi_6 <= 1'b0;
      state_0_6_lpi_6 <= 1'b0;
      state_0_7_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_4_lpi_6 <= 1'b0;
      state_0_5_lpi_6 <= 1'b0;
      state_0_6_lpi_6 <= 1'b0;
      state_0_7_lpi_6 <= 1'b0;
    end
    else if ( state_and_4_cse ) begin
      state_0_4_lpi_6 <= mux1h_4_nl & (~ (fsm_output[0]));
      state_0_5_lpi_6 <= mux1h_5_nl & (~ (fsm_output[0]));
      state_0_6_lpi_6 <= mux1h_6_nl & (~ (fsm_output[0]));
      state_0_7_lpi_6 <= mux1h_7_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_2_10_1_lpi_4 <= 1'b0;
      state_2_11_1_lpi_4 <= 1'b0;
      state_2_12_1_lpi_4 <= 1'b0;
      state_2_13_1_lpi_4 <= 1'b0;
      state_2_14_1_lpi_4 <= 1'b0;
      state_2_15_1_lpi_4 <= 1'b0;
      state_2_16_1_lpi_4 <= 1'b0;
      state_2_17_1_lpi_4 <= 1'b0;
      state_2_18_1_lpi_4 <= 1'b0;
      state_2_19_1_lpi_4 <= 1'b0;
      state_2_20_1_lpi_4 <= 1'b0;
      state_2_21_1_lpi_4 <= 1'b0;
      state_2_22_1_lpi_4 <= 1'b0;
      state_2_23_1_lpi_4 <= 1'b0;
      state_2_24_1_lpi_4 <= 1'b0;
      state_2_25_1_lpi_4 <= 1'b0;
    end
    else if ( rst ) begin
      state_2_10_1_lpi_4 <= 1'b0;
      state_2_11_1_lpi_4 <= 1'b0;
      state_2_12_1_lpi_4 <= 1'b0;
      state_2_13_1_lpi_4 <= 1'b0;
      state_2_14_1_lpi_4 <= 1'b0;
      state_2_15_1_lpi_4 <= 1'b0;
      state_2_16_1_lpi_4 <= 1'b0;
      state_2_17_1_lpi_4 <= 1'b0;
      state_2_18_1_lpi_4 <= 1'b0;
      state_2_19_1_lpi_4 <= 1'b0;
      state_2_20_1_lpi_4 <= 1'b0;
      state_2_21_1_lpi_4 <= 1'b0;
      state_2_22_1_lpi_4 <= 1'b0;
      state_2_23_1_lpi_4 <= 1'b0;
      state_2_24_1_lpi_4 <= 1'b0;
      state_2_25_1_lpi_4 <= 1'b0;
    end
    else if ( state_and_8_cse ) begin
      state_2_10_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[10]), state_xnor_nl, state_xnor_1_nl,
          xor_53_nl, state_4_16_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_11_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[11]), state_xnor_2_nl, state_xnor_3_nl,
          xor_51_nl, state_4_17_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_12_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[12]), state_xnor_4_nl, state_xnor_5_nl,
          xor_49_nl, state_4_18_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_13_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[13]), state_xnor_6_nl, state_xnor_7_nl,
          xor_47_nl, state_4_19_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_14_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[14]), state_xnor_8_nl, state_xnor_9_nl,
          xor_45_nl, state_4_2_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_15_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[15]), state_xnor_10_nl, state_xnor_11_nl,
          xor_43_nl, state_4_20_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_16_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[16]), state_xnor_12_nl, state_xnor_13_nl,
          xor_41_nl, state_4_21_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_17_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[17]), state_xnor_14_nl, state_xnor_15_nl,
          xor_39_nl, state_4_22_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_18_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[18]), state_xnor_16_nl, state_xnor_17_nl,
          xor_37_nl, state_4_4_23_sva_1_mx0w4, {(fsm_output[0]) , (fsm_output[1])
          , or_tmp_382 , and_885_cse , and_94_cse});
      state_2_19_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[19]), state_xnor_18_nl, state_xnor_19_nl,
          xor_35_nl, state_4_4_24_sva_1_mx0w4, {(fsm_output[0]) , (fsm_output[1])
          , or_tmp_382 , and_885_cse , and_94_cse});
      state_2_20_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[20]), state_xnor_20_nl, state_xnor_21_nl,
          xor_33_nl, state_4_25_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_21_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[21]), state_xnor_22_nl, state_xnor_23_nl,
          xor_31_nl, state_4_26_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_22_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[22]), state_xnor_24_nl, state_xnor_25_nl,
          xor_29_nl, state_4_27_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_23_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[23]), state_xnor_26_nl, state_xnor_27_nl,
          xor_27_nl, state_4_28_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_24_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[24]), state_xnor_28_nl, state_xnor_29_nl,
          xor_25_nl, state_4_29_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
      state_2_25_1_lpi_4 <= MUX1HOT_s_1_5_2((key4[25]), state_xnor_30_nl, state_xnor_31_nl,
          xor_23_nl, state_4_3_sva_2_mx0w4, {(fsm_output[0]) , (fsm_output[1]) ,
          or_tmp_382 , and_885_cse , and_94_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_2_26_1_lpi_4 <= 1'b0;
      state_2_27_1_lpi_4 <= 1'b0;
      state_2_28_1_lpi_4 <= 1'b0;
      state_2_29_1_lpi_4 <= 1'b0;
      state_2_30_1_lpi_4 <= 1'b0;
      state_2_31_1_lpi_4 <= 1'b0;
      state_2_32_1_lpi_4 <= 1'b0;
      state_2_33_1_lpi_4 <= 1'b0;
      state_2_34_1_lpi_4 <= 1'b0;
      state_2_35_1_lpi_4 <= 1'b0;
      state_2_36_1_lpi_4 <= 1'b0;
      state_2_37_1_lpi_4 <= 1'b0;
      state_2_38_1_lpi_4 <= 1'b0;
      state_2_39_1_lpi_4 <= 1'b0;
      state_2_40_1_lpi_4 <= 1'b0;
      state_2_41_1_lpi_4 <= 1'b0;
      state_2_42_1_lpi_4 <= 1'b0;
      state_2_43_1_lpi_4 <= 1'b0;
      state_2_44_1_lpi_4 <= 1'b0;
      state_2_45_1_lpi_4 <= 1'b0;
      state_2_46_1_lpi_4 <= 1'b0;
      state_2_47_1_lpi_4 <= 1'b0;
      state_2_48_1_lpi_4 <= 1'b0;
      state_2_49_1_lpi_4 <= 1'b0;
      state_2_50_1_lpi_4 <= 1'b0;
      state_2_51_1_lpi_4 <= 1'b0;
      state_2_52_1_lpi_4 <= 1'b0;
      state_2_53_1_lpi_4 <= 1'b0;
      state_2_54_1_lpi_4 <= 1'b0;
      state_2_55_1_lpi_4 <= 1'b0;
      state_2_56_1_lpi_4 <= 1'b0;
      state_2_57_1_lpi_4 <= 1'b0;
      state_2_8_1_lpi_4 <= 1'b0;
      state_2_9_1_lpi_4 <= 1'b0;
    end
    else if ( rst ) begin
      state_2_26_1_lpi_4 <= 1'b0;
      state_2_27_1_lpi_4 <= 1'b0;
      state_2_28_1_lpi_4 <= 1'b0;
      state_2_29_1_lpi_4 <= 1'b0;
      state_2_30_1_lpi_4 <= 1'b0;
      state_2_31_1_lpi_4 <= 1'b0;
      state_2_32_1_lpi_4 <= 1'b0;
      state_2_33_1_lpi_4 <= 1'b0;
      state_2_34_1_lpi_4 <= 1'b0;
      state_2_35_1_lpi_4 <= 1'b0;
      state_2_36_1_lpi_4 <= 1'b0;
      state_2_37_1_lpi_4 <= 1'b0;
      state_2_38_1_lpi_4 <= 1'b0;
      state_2_39_1_lpi_4 <= 1'b0;
      state_2_40_1_lpi_4 <= 1'b0;
      state_2_41_1_lpi_4 <= 1'b0;
      state_2_42_1_lpi_4 <= 1'b0;
      state_2_43_1_lpi_4 <= 1'b0;
      state_2_44_1_lpi_4 <= 1'b0;
      state_2_45_1_lpi_4 <= 1'b0;
      state_2_46_1_lpi_4 <= 1'b0;
      state_2_47_1_lpi_4 <= 1'b0;
      state_2_48_1_lpi_4 <= 1'b0;
      state_2_49_1_lpi_4 <= 1'b0;
      state_2_50_1_lpi_4 <= 1'b0;
      state_2_51_1_lpi_4 <= 1'b0;
      state_2_52_1_lpi_4 <= 1'b0;
      state_2_53_1_lpi_4 <= 1'b0;
      state_2_54_1_lpi_4 <= 1'b0;
      state_2_55_1_lpi_4 <= 1'b0;
      state_2_56_1_lpi_4 <= 1'b0;
      state_2_57_1_lpi_4 <= 1'b0;
      state_2_8_1_lpi_4 <= 1'b0;
      state_2_9_1_lpi_4 <= 1'b0;
    end
    else if ( state_and_24_cse ) begin
      state_2_26_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[26]), state_xnor_32_nl, state_xnor_33_nl,
          xor_21_nl, state_xnor_34_nl, state_4_30_sva_2_mx0w5, {(fsm_output[0]) ,
          (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_27_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[27]), state_xnor_35_nl, state_xnor_36_nl,
          xor_19_nl, state_xnor_37_nl, state_4_31_sva_2_mx0w5, {(fsm_output[0]) ,
          (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_28_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[28]), state_xnor_38_nl, state_xnor_39_nl,
          xor_17_nl, state_xnor_40_nl, state_4_4_sva_2_mx0w5, {(fsm_output[0]) ,
          (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_29_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[29]), state_xnor_41_nl, state_xnor_42_nl,
          xor_15_nl, state_xnor_43_nl, state_4_5_sva_2_mx0w5, {(fsm_output[0]) ,
          (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_30_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[30]), state_xnor_44_nl, state_xnor_45_nl,
          xor_13_nl, state_xnor_46_nl, state_4_6_sva_2_mx0w5, {(fsm_output[0]) ,
          (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_31_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[31]), state_xnor_47_nl, state_xnor_48_nl,
          xor_7_nl, state_xnor_49_nl, state_4_7_sva_2_mx0w5, {(fsm_output[0]) , (fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_32_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[0]), state_xnor_50_nl, state_xnor_51_nl,
          data_out_rsci_idat_0_mx0w6, state_xnor_52_nl, state_4_32_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_33_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[1]), state_xnor_53_nl, state_xnor_54_nl,
          data_out_rsci_idat_1_mx0w6, state_xnor_55_nl, state_4_33_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_34_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[2]), state_xnor_56_nl, state_xnor_57_nl,
          data_out_rsci_idat_2_mx0w6, state_xnor_58_nl, state_4_34_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_35_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[3]), state_xnor_59_nl, state_xnor_60_nl,
          data_out_rsci_idat_3_mx0w6, state_xnor_61_nl, state_4_35_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_36_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[4]), state_xnor_62_nl, state_xnor_63_nl,
          data_out_rsci_idat_4_mx0w6, state_xnor_64_nl, state_4_36_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_37_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[5]), state_xnor_65_nl, state_xnor_66_nl,
          data_out_rsci_idat_5_mx0w6, state_xnor_67_nl, state_4_37_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_38_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[6]), state_xnor_68_nl, state_xnor_69_nl,
          data_out_rsci_idat_6_mx0w6, state_xnor_70_nl, state_4_38_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_39_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[7]), state_xnor_71_nl, state_xnor_72_nl,
          data_out_rsci_idat_7_mx0w6, state_xnor_73_nl, state_4_39_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_40_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[8]), state_xnor_74_nl, state_xnor_75_nl,
          data_out_rsci_idat_8_mx0w6, state_xnor_76_nl, state_4_40_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_41_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[9]), state_xnor_77_nl, state_xnor_78_nl,
          data_out_rsci_idat_9_mx0w6, state_xnor_79_nl, state_4_41_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_42_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[10]), state_xnor_80_nl, state_xnor_81_nl,
          data_out_rsci_idat_10_mx0w6, state_xnor_82_nl, state_4_42_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_43_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[11]), state_xnor_83_nl, state_xnor_84_nl,
          data_out_rsci_idat_11_mx0w6, state_xnor_85_nl, state_4_43_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_44_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[12]), state_xnor_86_nl, state_xnor_87_nl,
          data_out_rsci_idat_12_mx0w6, state_xnor_88_nl, state_4_44_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_45_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[13]), state_xnor_89_nl, state_xnor_90_nl,
          data_out_rsci_idat_13_mx0w6, state_xnor_91_nl, state_4_45_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_46_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[14]), state_xnor_92_nl, state_xnor_93_nl,
          data_out_rsci_idat_14_mx0w6, state_xnor_94_nl, state_4_46_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_47_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[15]), state_xnor_95_nl, state_xnor_96_nl,
          data_out_rsci_idat_15_mx0w6, state_xnor_97_nl, state_4_47_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_48_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[16]), state_xnor_98_nl, state_xnor_99_nl,
          data_out_rsci_idat_16_mx0w6, state_xnor_100_nl, state_4_48_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_49_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[17]), state_xnor_101_nl, state_xnor_102_nl,
          data_out_rsci_idat_17_mx0w6, state_xnor_103_nl, state_4_49_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_50_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[18]), state_xnor_104_nl, state_xnor_105_nl,
          data_out_rsci_idat_18_mx0w6, state_xnor_106_nl, state_4_50_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_51_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[19]), state_xnor_107_nl, state_xnor_108_nl,
          data_out_rsci_idat_19_mx0w6, state_xnor_109_nl, state_4_51_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_52_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[20]), state_xnor_110_nl, state_xnor_111_nl,
          data_out_rsci_idat_20_mx0w6, state_xnor_112_nl, state_4_52_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_53_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[21]), state_xnor_113_nl, state_xnor_114_nl,
          data_out_rsci_idat_21_mx0w6, state_xnor_115_nl, state_4_53_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_54_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[22]), state_xnor_116_nl, state_xnor_117_nl,
          data_out_rsci_idat_22_mx0w6, state_xnor_118_nl, state_4_54_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_55_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[23]), state_xnor_119_nl, state_xnor_120_nl,
          data_out_rsci_idat_23_mx0w6, state_xnor_121_nl, state_4_55_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_56_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[24]), state_xnor_122_nl, state_xnor_123_nl,
          data_out_rsci_idat_24_mx0w6, state_xnor_124_nl, state_4_56_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_57_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[25]), state_xnor_125_nl, state_xnor_126_nl,
          data_out_rsci_idat_25_mx0w6, state_xnor_127_nl, state_4_57_sva_2_mx0w5,
          {(fsm_output[0]) , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse
          , and_94_cse});
      state_2_8_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[8]), state_xnor_146_nl, state_xnor_147_nl,
          data_out_rsci_idat_8_mx0w7, state_xnor_148_nl, state_4_8_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_2_9_1_lpi_4 <= MUX1HOT_s_1_6_2((key4[9]), state_xnor_149_nl, state_xnor_150_nl,
          data_out_rsci_idat_9_mx0w7, state_xnor_151_nl, state_4_9_sva_2_mx0w5, {(fsm_output[0])
          , (fsm_output[1]) , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_2_58_1_lpi_4 <= 1'b0;
      state_2_59_1_lpi_4 <= 1'b0;
      state_2_60_1_lpi_4 <= 1'b0;
      state_2_61_1_lpi_4 <= 1'b0;
      state_2_62_1_lpi_4 <= 1'b0;
      state_2_63_1_lpi_4 <= 1'b0;
    end
    else if ( rst ) begin
      state_2_58_1_lpi_4 <= 1'b0;
      state_2_59_1_lpi_4 <= 1'b0;
      state_2_60_1_lpi_4 <= 1'b0;
      state_2_61_1_lpi_4 <= 1'b0;
      state_2_62_1_lpi_4 <= 1'b0;
      state_2_63_1_lpi_4 <= 1'b0;
    end
    else if ( state_and_56_cse ) begin
      state_2_58_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[26]), state_xnor_128_nl, state_xnor_129_nl,
          Encrypt_Top_linear_2_xnor_nl, xor_64_nl, state_xnor_130_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
      state_2_59_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[27]), state_xnor_131_nl, state_xnor_132_nl,
          Encrypt_Top_linear_2_xnor_1_nl, xor_66_nl, state_xnor_133_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
      state_2_60_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[28]), state_xnor_134_nl, state_xnor_135_nl,
          Encrypt_Top_linear_2_xnor_2_nl, xor_68_nl, state_xnor_136_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
      state_2_61_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[29]), state_xnor_137_nl, state_xnor_138_nl,
          Encrypt_Top_linear_2_xnor_3_nl, xor_70_nl, state_xnor_139_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
      state_2_62_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[30]), state_xnor_140_nl, state_xnor_141_nl,
          Encrypt_Top_linear_2_xnor_4_nl, xor_72_nl, state_xnor_142_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
      state_2_63_1_lpi_4 <= MUX1HOT_s_1_6_2((key3[31]), state_xnor_143_nl, state_xnor_144_nl,
          Encrypt_Top_linear_2_xnor_5_nl, xor_74_nl, state_xnor_145_nl, {(fsm_output[0])
          , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse ,
          (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_10_lpi_6 <= 1'b0;
      state_0_11_lpi_6 <= 1'b0;
      state_0_12_lpi_6 <= 1'b0;
      state_0_13_lpi_6 <= 1'b0;
      state_0_14_lpi_6 <= 1'b0;
      state_0_15_lpi_6 <= 1'b0;
      state_0_16_lpi_6 <= 1'b0;
      state_0_17_lpi_6 <= 1'b0;
      state_0_18_lpi_6 <= 1'b0;
      state_0_19_lpi_6 <= 1'b0;
      state_0_20_lpi_6 <= 1'b0;
      state_0_21_lpi_6 <= 1'b0;
      state_0_22_lpi_6 <= 1'b0;
      state_0_23_lpi_6 <= 1'b0;
      state_0_24_lpi_6 <= 1'b0;
      state_0_25_lpi_6 <= 1'b0;
      state_0_26_lpi_6 <= 1'b0;
      state_0_27_lpi_6 <= 1'b0;
      state_0_28_lpi_6 <= 1'b0;
      state_0_29_lpi_6 <= 1'b0;
      state_0_30_lpi_6 <= 1'b0;
      state_0_31_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_10_lpi_6 <= 1'b0;
      state_0_11_lpi_6 <= 1'b0;
      state_0_12_lpi_6 <= 1'b0;
      state_0_13_lpi_6 <= 1'b0;
      state_0_14_lpi_6 <= 1'b0;
      state_0_15_lpi_6 <= 1'b0;
      state_0_16_lpi_6 <= 1'b0;
      state_0_17_lpi_6 <= 1'b0;
      state_0_18_lpi_6 <= 1'b0;
      state_0_19_lpi_6 <= 1'b0;
      state_0_20_lpi_6 <= 1'b0;
      state_0_21_lpi_6 <= 1'b0;
      state_0_22_lpi_6 <= 1'b0;
      state_0_23_lpi_6 <= 1'b0;
      state_0_24_lpi_6 <= 1'b0;
      state_0_25_lpi_6 <= 1'b0;
      state_0_26_lpi_6 <= 1'b0;
      state_0_27_lpi_6 <= 1'b0;
      state_0_28_lpi_6 <= 1'b0;
      state_0_29_lpi_6 <= 1'b0;
      state_0_30_lpi_6 <= 1'b0;
      state_0_31_lpi_6 <= 1'b0;
    end
    else if ( state_and_64_cse ) begin
      state_0_10_lpi_6 <= mux1h_64_nl & (~ (fsm_output[0]));
      state_0_11_lpi_6 <= mux1h_65_nl & (~ (fsm_output[0]));
      state_0_12_lpi_6 <= mux1h_66_nl & (~ (fsm_output[0]));
      state_0_13_lpi_6 <= mux1h_67_nl & (~ (fsm_output[0]));
      state_0_14_lpi_6 <= mux1h_68_nl & (~ (fsm_output[0]));
      state_0_15_lpi_6 <= mux1h_69_nl & (~ (fsm_output[0]));
      state_0_16_lpi_6 <= mux1h_70_nl & (~ (fsm_output[0]));
      state_0_17_lpi_6 <= mux1h_71_nl & (~ (fsm_output[0]));
      state_0_18_lpi_6 <= mux1h_72_nl & (~ (fsm_output[0]));
      state_0_19_lpi_6 <= mux1h_73_nl & (~ (fsm_output[0]));
      state_0_20_lpi_6 <= mux1h_74_nl & (~ (fsm_output[0]));
      state_0_21_lpi_6 <= mux1h_75_nl & (~ (fsm_output[0]));
      state_0_22_lpi_6 <= mux1h_76_nl & (~ (fsm_output[0]));
      state_0_23_lpi_6 <= mux1h_77_nl & (~ (fsm_output[0]));
      state_0_24_lpi_6 <= mux1h_78_nl & (~ (fsm_output[0]));
      state_0_25_lpi_6 <= mux1h_79_nl & (~ (fsm_output[0]));
      state_0_26_lpi_6 <= mux1h_80_nl & (~ (fsm_output[0]));
      state_0_27_lpi_6 <= mux1h_81_nl & (~ (fsm_output[0]));
      state_0_28_lpi_6 <= mux1h_82_nl & (~ (fsm_output[0]));
      state_0_29_lpi_6 <= mux1h_83_nl & (~ (fsm_output[0]));
      state_0_30_lpi_6 <= mux1h_84_nl & (~ (fsm_output[0]));
      state_0_31_lpi_6 <= mux1h_85_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_32_lpi_6 <= 1'b0;
      state_0_33_lpi_6 <= 1'b0;
      state_0_34_lpi_6 <= 1'b0;
      state_0_35_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_32_lpi_6 <= 1'b0;
      state_0_33_lpi_6 <= 1'b0;
      state_0_34_lpi_6 <= 1'b0;
      state_0_35_lpi_6 <= 1'b0;
    end
    else if ( state_and_86_cse ) begin
      state_0_32_lpi_6 <= mux1h_86_nl & (~ (fsm_output[0]));
      state_0_33_lpi_6 <= mux1h_87_nl | (fsm_output[0]);
      state_0_34_lpi_6 <= mux1h_88_nl | (fsm_output[0]);
      state_0_35_lpi_6 <= mux1h_89_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_36_lpi_6 <= 1'b0;
      state_0_37_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_36_lpi_6 <= 1'b0;
      state_0_37_lpi_6 <= 1'b0;
    end
    else if ( state_and_90_cse ) begin
      state_0_36_lpi_6 <= mux1h_90_nl & (~ (fsm_output[0]));
      state_0_37_lpi_6 <= mux1h_91_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_38_lpi_6 <= 1'b0;
      state_0_39_lpi_6 <= 1'b0;
      state_0_40_lpi_6 <= 1'b0;
      state_0_41_lpi_6 <= 1'b0;
      state_0_42_lpi_6 <= 1'b0;
      state_0_43_lpi_6 <= 1'b0;
      state_0_45_lpi_6 <= 1'b0;
      state_0_46_lpi_6 <= 1'b0;
      state_0_47_lpi_6 <= 1'b0;
      state_0_48_lpi_6 <= 1'b0;
      state_0_49_lpi_6 <= 1'b0;
      state_0_50_lpi_6 <= 1'b0;
      state_0_51_lpi_6 <= 1'b0;
      state_0_52_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_38_lpi_6 <= 1'b0;
      state_0_39_lpi_6 <= 1'b0;
      state_0_40_lpi_6 <= 1'b0;
      state_0_41_lpi_6 <= 1'b0;
      state_0_42_lpi_6 <= 1'b0;
      state_0_43_lpi_6 <= 1'b0;
      state_0_45_lpi_6 <= 1'b0;
      state_0_46_lpi_6 <= 1'b0;
      state_0_47_lpi_6 <= 1'b0;
      state_0_48_lpi_6 <= 1'b0;
      state_0_49_lpi_6 <= 1'b0;
      state_0_50_lpi_6 <= 1'b0;
      state_0_51_lpi_6 <= 1'b0;
      state_0_52_lpi_6 <= 1'b0;
    end
    else if ( state_and_92_cse ) begin
      state_0_38_lpi_6 <= mux1h_92_nl & (~ (fsm_output[0]));
      state_0_39_lpi_6 <= mux1h_93_nl & (~ (fsm_output[0]));
      state_0_40_lpi_6 <= mux1h_94_nl & (~ (fsm_output[0]));
      state_0_41_lpi_6 <= mux1h_95_nl & (~ (fsm_output[0]));
      state_0_42_lpi_6 <= mux1h_96_nl | (fsm_output[0]);
      state_0_43_lpi_6 <= mux1h_97_nl | (fsm_output[0]);
      state_0_45_lpi_6 <= mux1h_99_nl & (~ (fsm_output[0]));
      state_0_46_lpi_6 <= mux1h_100_nl & (~ (fsm_output[0]));
      state_0_47_lpi_6 <= mux1h_101_nl & (~ (fsm_output[0]));
      state_0_48_lpi_6 <= mux1h_102_nl & (~ (fsm_output[0]));
      state_0_49_lpi_6 <= mux1h_103_nl & (~ (fsm_output[0]));
      state_0_50_lpi_6 <= mux1h_104_nl & (~ (fsm_output[0]));
      state_0_51_lpi_6 <= mux1h_105_nl & (~ (fsm_output[0]));
      state_0_52_lpi_6 <= mux1h_106_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_44_lpi_6 <= 1'b0;
      state_0_53_lpi_6 <= 1'b0;
      state_0_54_lpi_6 <= 1'b0;
      state_0_55_lpi_6 <= 1'b0;
      state_0_56_lpi_6 <= 1'b0;
      state_0_57_lpi_6 <= 1'b0;
      state_0_58_lpi_6 <= 1'b0;
      state_0_59_lpi_6 <= 1'b0;
      state_0_60_lpi_6 <= 1'b0;
      state_0_61_lpi_6 <= 1'b0;
      state_0_62_lpi_6 <= 1'b0;
      state_0_63_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_44_lpi_6 <= 1'b0;
      state_0_53_lpi_6 <= 1'b0;
      state_0_54_lpi_6 <= 1'b0;
      state_0_55_lpi_6 <= 1'b0;
      state_0_56_lpi_6 <= 1'b0;
      state_0_57_lpi_6 <= 1'b0;
      state_0_58_lpi_6 <= 1'b0;
      state_0_59_lpi_6 <= 1'b0;
      state_0_60_lpi_6 <= 1'b0;
      state_0_61_lpi_6 <= 1'b0;
      state_0_62_lpi_6 <= 1'b0;
      state_0_63_lpi_6 <= 1'b0;
    end
    else if ( state_and_98_cse ) begin
      state_0_44_lpi_6 <= mux1h_98_nl & (~ (fsm_output[0]));
      state_0_53_lpi_6 <= mux1h_107_nl & (~ (fsm_output[0]));
      state_0_54_lpi_6 <= mux1h_108_nl | (fsm_output[0]);
      state_0_55_lpi_6 <= mux1h_109_nl & (~ (fsm_output[0]));
      state_0_56_lpi_6 <= mux1h_110_nl & (~ (fsm_output[0]));
      state_0_57_lpi_6 <= mux1h_111_nl & (~ (fsm_output[0]));
      state_0_58_lpi_6 <= mux1h_112_nl & (~ (fsm_output[0]));
      state_0_59_lpi_6 <= mux1h_113_nl & (~ (fsm_output[0]));
      state_0_60_lpi_6 <= mux1h_114_nl & (~ (fsm_output[0]));
      state_0_61_lpi_6 <= mux1h_115_nl & (~ (fsm_output[0]));
      state_0_62_lpi_6 <= mux1h_116_nl & (~ (fsm_output[0]));
      state_0_63_lpi_6 <= mux1h_117_nl | (fsm_output[0]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_0_8_lpi_6 <= 1'b0;
      state_0_9_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_0_8_lpi_6 <= 1'b0;
      state_0_9_lpi_6 <= 1'b0;
    end
    else if ( state_and_118_cse ) begin
      state_0_8_lpi_6 <= mux1h_118_nl & (~ (fsm_output[0]));
      state_0_9_lpi_6 <= mux1h_119_nl & (~ (fsm_output[0]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_2_0_1_lpi_4 <= 1'b0;
      state_2_1_1_lpi_4 <= 1'b0;
      state_2_2_1_lpi_4 <= 1'b0;
      state_2_3_1_lpi_4 <= 1'b0;
      state_2_4_1_lpi_4 <= 1'b0;
      state_2_5_1_lpi_4 <= 1'b0;
      state_2_6_1_lpi_4 <= 1'b0;
      state_2_7_1_lpi_4 <= 1'b0;
    end
    else if ( rst ) begin
      state_2_0_1_lpi_4 <= 1'b0;
      state_2_1_1_lpi_4 <= 1'b0;
      state_2_2_1_lpi_4 <= 1'b0;
      state_2_3_1_lpi_4 <= 1'b0;
      state_2_4_1_lpi_4 <= 1'b0;
      state_2_5_1_lpi_4 <= 1'b0;
      state_2_6_1_lpi_4 <= 1'b0;
      state_2_7_1_lpi_4 <= 1'b0;
    end
    else if ( state_and_120_cse ) begin
      state_2_0_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[0]), state_xnor_152_nl, state_2_0_1_sva_4,
          state_2_0_1_lpi_6, data_out_rsci_idat_0_mx0w7, state_xnor_153_nl, state_3_0_sva_3_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_1_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[1]), state_xnor_155_nl, state_2_1_1_sva_4,
          state_2_1_1_lpi_6, data_out_rsci_idat_1_mx0w7, state_xnor_156_nl, state_3_1_sva_3_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_2_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[2]), state_xnor_158_nl, state_2_2_1_sva_4,
          state_2_2_1_lpi_6, xor_69_nl, state_xnor_159_nl, state_3_10_sva_2_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_3_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[3]), state_xnor_161_nl, state_2_3_1_sva_4,
          state_2_3_1_lpi_6, xor_67_nl, state_xnor_162_nl, state_3_11_sva_2_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_4_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[4]), state_xnor_164_nl, state_2_4_1_sva_4,
          state_2_4_1_lpi_6, xor_65_nl, state_xnor_165_nl, state_3_12_sva_2_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_5_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[5]), state_xnor_167_nl, state_2_5_1_sva_4,
          state_2_5_1_lpi_6, xor_63_nl, state_xnor_168_nl, state_3_13_sva_2_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_6_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[6]), state_xnor_170_nl, state_2_6_1_sva_4,
          state_2_6_1_lpi_6, xor_61_nl, state_xnor_171_nl, state_3_14_sva_2_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
      state_2_7_1_lpi_4 <= MUX1HOT_s_1_7_2((key4[7]), state_xnor_173_nl, state_2_7_1_sva_4,
          state_2_7_1_lpi_6, xor_59_nl, state_xnor_174_nl, state_3_15_sva_3_mx0w6,
          {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[4]) , (fsm_output[5])
          , (fsm_output[13]) , and_39_cse , and_94_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      plaintext_31_0_sva_31 <= 1'b0;
      plaintext_31_0_sva_30 <= 1'b0;
      plaintext_31_0_sva_29 <= 1'b0;
      plaintext_31_0_sva_28 <= 1'b0;
      plaintext_31_0_sva_27 <= 1'b0;
      plaintext_31_0_sva_26 <= 1'b0;
      plaintext_31_0_sva_25 <= 1'b0;
      plaintext_31_0_sva_24 <= 1'b0;
      plaintext_31_0_sva_23 <= 1'b0;
      plaintext_31_0_sva_22 <= 1'b0;
      plaintext_31_0_sva_21 <= 1'b0;
      plaintext_31_0_sva_20 <= 1'b0;
      plaintext_31_0_sva_19 <= 1'b0;
      plaintext_31_0_sva_18 <= 1'b0;
      plaintext_31_0_sva_17 <= 1'b0;
      plaintext_31_0_sva_16 <= 1'b0;
      plaintext_31_0_sva_15 <= 1'b0;
      plaintext_31_0_sva_14 <= 1'b0;
      plaintext_31_0_sva_13 <= 1'b0;
      plaintext_31_0_sva_12 <= 1'b0;
      plaintext_31_0_sva_11 <= 1'b0;
      plaintext_31_0_sva_10 <= 1'b0;
      plaintext_31_0_sva_9 <= 1'b0;
      plaintext_31_0_sva_8 <= 1'b0;
      plaintext_31_0_sva_7 <= 1'b0;
      plaintext_31_0_sva_6 <= 1'b0;
      plaintext_31_0_sva_5 <= 1'b0;
      plaintext_31_0_sva_4 <= 1'b0;
      plaintext_31_0_sva_3 <= 1'b0;
      plaintext_31_0_sva_2 <= 1'b0;
      plaintext_31_0_sva_1 <= 1'b0;
      plaintext_31_0_sva_0 <= 1'b0;
    end
    else if ( rst ) begin
      plaintext_31_0_sva_31 <= 1'b0;
      plaintext_31_0_sva_30 <= 1'b0;
      plaintext_31_0_sva_29 <= 1'b0;
      plaintext_31_0_sva_28 <= 1'b0;
      plaintext_31_0_sva_27 <= 1'b0;
      plaintext_31_0_sva_26 <= 1'b0;
      plaintext_31_0_sva_25 <= 1'b0;
      plaintext_31_0_sva_24 <= 1'b0;
      plaintext_31_0_sva_23 <= 1'b0;
      plaintext_31_0_sva_22 <= 1'b0;
      plaintext_31_0_sva_21 <= 1'b0;
      plaintext_31_0_sva_20 <= 1'b0;
      plaintext_31_0_sva_19 <= 1'b0;
      plaintext_31_0_sva_18 <= 1'b0;
      plaintext_31_0_sva_17 <= 1'b0;
      plaintext_31_0_sva_16 <= 1'b0;
      plaintext_31_0_sva_15 <= 1'b0;
      plaintext_31_0_sva_14 <= 1'b0;
      plaintext_31_0_sva_13 <= 1'b0;
      plaintext_31_0_sva_12 <= 1'b0;
      plaintext_31_0_sva_11 <= 1'b0;
      plaintext_31_0_sva_10 <= 1'b0;
      plaintext_31_0_sva_9 <= 1'b0;
      plaintext_31_0_sva_8 <= 1'b0;
      plaintext_31_0_sva_7 <= 1'b0;
      plaintext_31_0_sva_6 <= 1'b0;
      plaintext_31_0_sva_5 <= 1'b0;
      plaintext_31_0_sva_4 <= 1'b0;
      plaintext_31_0_sva_3 <= 1'b0;
      plaintext_31_0_sva_2 <= 1'b0;
      plaintext_31_0_sva_1 <= 1'b0;
      plaintext_31_0_sva_0 <= 1'b0;
    end
    else if ( plaintext_and_ssc ) begin
      plaintext_31_0_sva_31 <= MUX1HOT_s_1_3_2((key2[31]), state_1_1_31_0_sva_1_31_1,
          (data_in_rsci_idat_mxwt[31]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_30 <= MUX1HOT_s_1_3_2((key2[30]), state_1_1_31_0_sva_1_30_1,
          (data_in_rsci_idat_mxwt[30]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_29 <= MUX1HOT_s_1_3_2((key2[29]), state_1_1_31_0_sva_1_29_1,
          (data_in_rsci_idat_mxwt[29]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_28 <= MUX1HOT_s_1_3_2((key2[28]), state_1_1_31_0_sva_1_28_1,
          (data_in_rsci_idat_mxwt[28]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_27 <= MUX1HOT_s_1_3_2((key2[27]), state_1_1_31_0_sva_1_27_1,
          (data_in_rsci_idat_mxwt[27]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_26 <= MUX1HOT_s_1_3_2((key2[26]), state_1_1_31_0_sva_1_26_1,
          (data_in_rsci_idat_mxwt[26]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_25 <= MUX1HOT_s_1_3_2((key2[25]), state_1_1_31_0_sva_1_25_1,
          (data_in_rsci_idat_mxwt[25]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_24 <= MUX1HOT_s_1_3_2((key2[24]), state_1_1_31_0_sva_1_24_1,
          (data_in_rsci_idat_mxwt[24]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_23 <= MUX1HOT_s_1_3_2((key2[23]), state_1_1_31_0_sva_1_23_1,
          (data_in_rsci_idat_mxwt[23]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_22 <= MUX1HOT_s_1_3_2((key2[22]), state_1_1_31_0_sva_1_22_1,
          (data_in_rsci_idat_mxwt[22]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_21 <= MUX1HOT_s_1_3_2((key2[21]), state_1_1_31_0_sva_1_21_1,
          (data_in_rsci_idat_mxwt[21]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_20 <= MUX1HOT_s_1_3_2((key2[20]), state_1_1_31_0_sva_1_20_1,
          (data_in_rsci_idat_mxwt[20]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_19 <= MUX1HOT_s_1_3_2((key2[19]), state_1_1_31_0_sva_1_19_1,
          (data_in_rsci_idat_mxwt[19]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_18 <= MUX1HOT_s_1_3_2((key2[18]), state_1_1_31_0_sva_1_18_1,
          (data_in_rsci_idat_mxwt[18]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_17 <= MUX1HOT_s_1_3_2((key2[17]), state_1_1_31_0_sva_1_17_1,
          (data_in_rsci_idat_mxwt[17]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_16 <= MUX1HOT_s_1_3_2((key2[16]), state_1_1_31_0_sva_1_16_1,
          (data_in_rsci_idat_mxwt[16]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_15 <= MUX1HOT_s_1_3_2((key2[15]), state_1_1_31_0_sva_1_15_1,
          (data_in_rsci_idat_mxwt[15]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_14 <= MUX1HOT_s_1_3_2((key2[14]), state_1_1_31_0_sva_1_14_1,
          (data_in_rsci_idat_mxwt[14]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_13 <= MUX1HOT_s_1_3_2((key2[13]), state_1_1_31_0_sva_1_13_1,
          (data_in_rsci_idat_mxwt[13]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_12 <= MUX1HOT_s_1_3_2((key2[12]), state_1_1_31_0_sva_1_12_1,
          (data_in_rsci_idat_mxwt[12]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_11 <= MUX1HOT_s_1_3_2((key2[11]), state_1_1_31_0_sva_1_11_1,
          (data_in_rsci_idat_mxwt[11]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_10 <= MUX1HOT_s_1_3_2((key2[10]), state_1_1_31_0_sva_1_10_1,
          (data_in_rsci_idat_mxwt[10]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_9 <= MUX1HOT_s_1_3_2((key2[9]), state_1_1_31_0_sva_1_9_1,
          (data_in_rsci_idat_mxwt[9]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_8 <= MUX1HOT_s_1_3_2((key2[8]), state_1_1_31_0_sva_1_8_1,
          (data_in_rsci_idat_mxwt[8]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_7 <= MUX1HOT_s_1_3_2((key2[7]), state_1_1_31_0_sva_1_7_1,
          (data_in_rsci_idat_mxwt[7]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_6 <= MUX1HOT_s_1_3_2((key2[6]), state_1_1_31_0_sva_1_6_1,
          (data_in_rsci_idat_mxwt[6]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_5 <= MUX1HOT_s_1_3_2((key2[5]), state_1_1_31_0_sva_1_5_1,
          (data_in_rsci_idat_mxwt[5]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_4 <= MUX1HOT_s_1_3_2((key2[4]), state_1_1_31_0_sva_1_4_1,
          (data_in_rsci_idat_mxwt[4]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_3 <= MUX1HOT_s_1_3_2((key2[3]), state_1_1_31_0_sva_1_3_1,
          (data_in_rsci_idat_mxwt[3]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_2 <= MUX1HOT_s_1_3_2((key2[2]), state_1_1_31_0_sva_1_2_1,
          (data_in_rsci_idat_mxwt[2]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_1 <= MUX1HOT_s_1_3_2((key2[1]), state_1_1_31_0_sva_1_1_1,
          (data_in_rsci_idat_mxwt[1]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
      plaintext_31_0_sva_0 <= MUX1HOT_s_1_3_2((key2[0]), state_1_1_31_0_sva_1_0_1,
          (data_in_rsci_idat_mxwt[0]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[10])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      plaintext_63_32_sva_31 <= 1'b0;
      plaintext_63_32_sva_30 <= 1'b0;
      plaintext_63_32_sva_29 <= 1'b0;
      plaintext_63_32_sva_28 <= 1'b0;
      plaintext_63_32_sva_27 <= 1'b0;
      plaintext_63_32_sva_26 <= 1'b0;
      plaintext_63_32_sva_25 <= 1'b0;
      plaintext_63_32_sva_24 <= 1'b0;
      plaintext_63_32_sva_23 <= 1'b0;
      plaintext_63_32_sva_22 <= 1'b0;
      plaintext_63_32_sva_21 <= 1'b0;
      plaintext_63_32_sva_20 <= 1'b0;
      plaintext_63_32_sva_19 <= 1'b0;
      plaintext_63_32_sva_18 <= 1'b0;
      plaintext_63_32_sva_17 <= 1'b0;
      plaintext_63_32_sva_16 <= 1'b0;
      plaintext_63_32_sva_15 <= 1'b0;
      plaintext_63_32_sva_14 <= 1'b0;
      plaintext_63_32_sva_13 <= 1'b0;
      plaintext_63_32_sva_12 <= 1'b0;
      plaintext_63_32_sva_11 <= 1'b0;
      plaintext_63_32_sva_10 <= 1'b0;
      plaintext_63_32_sva_9 <= 1'b0;
      plaintext_63_32_sva_8 <= 1'b0;
      plaintext_63_32_sva_7 <= 1'b0;
      plaintext_63_32_sva_6 <= 1'b0;
      plaintext_63_32_sva_5 <= 1'b0;
      plaintext_63_32_sva_4 <= 1'b0;
      plaintext_63_32_sva_3 <= 1'b0;
      plaintext_63_32_sva_2 <= 1'b0;
      plaintext_63_32_sva_1 <= 1'b0;
      plaintext_63_32_sva_0 <= 1'b0;
    end
    else if ( rst ) begin
      plaintext_63_32_sva_31 <= 1'b0;
      plaintext_63_32_sva_30 <= 1'b0;
      plaintext_63_32_sva_29 <= 1'b0;
      plaintext_63_32_sva_28 <= 1'b0;
      plaintext_63_32_sva_27 <= 1'b0;
      plaintext_63_32_sva_26 <= 1'b0;
      plaintext_63_32_sva_25 <= 1'b0;
      plaintext_63_32_sva_24 <= 1'b0;
      plaintext_63_32_sva_23 <= 1'b0;
      plaintext_63_32_sva_22 <= 1'b0;
      plaintext_63_32_sva_21 <= 1'b0;
      plaintext_63_32_sva_20 <= 1'b0;
      plaintext_63_32_sva_19 <= 1'b0;
      plaintext_63_32_sva_18 <= 1'b0;
      plaintext_63_32_sva_17 <= 1'b0;
      plaintext_63_32_sva_16 <= 1'b0;
      plaintext_63_32_sva_15 <= 1'b0;
      plaintext_63_32_sva_14 <= 1'b0;
      plaintext_63_32_sva_13 <= 1'b0;
      plaintext_63_32_sva_12 <= 1'b0;
      plaintext_63_32_sva_11 <= 1'b0;
      plaintext_63_32_sva_10 <= 1'b0;
      plaintext_63_32_sva_9 <= 1'b0;
      plaintext_63_32_sva_8 <= 1'b0;
      plaintext_63_32_sva_7 <= 1'b0;
      plaintext_63_32_sva_6 <= 1'b0;
      plaintext_63_32_sva_5 <= 1'b0;
      plaintext_63_32_sva_4 <= 1'b0;
      plaintext_63_32_sva_3 <= 1'b0;
      plaintext_63_32_sva_2 <= 1'b0;
      plaintext_63_32_sva_1 <= 1'b0;
      plaintext_63_32_sva_0 <= 1'b0;
    end
    else if ( plaintext_and_1_ssc ) begin
      plaintext_63_32_sva_31 <= MUX1HOT_s_1_3_2((key1[31]), state_1_1_63_32_sva_1_31_1,
          (data_in_rsci_idat_mxwt[31]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_30 <= MUX1HOT_s_1_3_2((key1[30]), state_1_1_63_32_sva_1_30_1,
          (data_in_rsci_idat_mxwt[30]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_29 <= MUX1HOT_s_1_3_2((key1[29]), state_1_1_63_32_sva_1_29_1,
          (data_in_rsci_idat_mxwt[29]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_28 <= MUX1HOT_s_1_3_2((key1[28]), state_1_1_63_32_sva_1_28_1,
          (data_in_rsci_idat_mxwt[28]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_27 <= MUX1HOT_s_1_3_2((key1[27]), state_1_1_63_32_sva_1_27_1,
          (data_in_rsci_idat_mxwt[27]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_26 <= MUX1HOT_s_1_3_2((key1[26]), state_1_1_63_32_sva_1_26_1,
          (data_in_rsci_idat_mxwt[26]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_25 <= MUX1HOT_s_1_3_2((key1[25]), state_1_1_63_32_sva_1_25_1,
          (data_in_rsci_idat_mxwt[25]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_24 <= MUX1HOT_s_1_3_2((key1[24]), state_1_1_63_32_sva_1_24_1,
          (data_in_rsci_idat_mxwt[24]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_23 <= MUX1HOT_s_1_3_2((key1[23]), state_1_1_63_32_sva_1_23_1,
          (data_in_rsci_idat_mxwt[23]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_22 <= MUX1HOT_s_1_3_2((key1[22]), state_1_1_63_32_sva_1_22_1,
          (data_in_rsci_idat_mxwt[22]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_21 <= MUX1HOT_s_1_3_2((key1[21]), state_1_1_63_32_sva_1_21_1,
          (data_in_rsci_idat_mxwt[21]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_20 <= MUX1HOT_s_1_3_2((key1[20]), state_1_1_63_32_sva_1_20_1,
          (data_in_rsci_idat_mxwt[20]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_19 <= MUX1HOT_s_1_3_2((key1[19]), state_1_1_63_32_sva_1_19_1,
          (data_in_rsci_idat_mxwt[19]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_18 <= MUX1HOT_s_1_3_2((key1[18]), state_1_1_63_32_sva_1_18_1,
          (data_in_rsci_idat_mxwt[18]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_17 <= MUX1HOT_s_1_3_2((key1[17]), state_1_1_63_32_sva_1_17_1,
          (data_in_rsci_idat_mxwt[17]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_16 <= MUX1HOT_s_1_3_2((key1[16]), state_1_1_63_32_sva_1_16_1,
          (data_in_rsci_idat_mxwt[16]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_15 <= MUX1HOT_s_1_3_2((key1[15]), state_1_1_63_32_sva_1_15_1,
          (data_in_rsci_idat_mxwt[15]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_14 <= MUX1HOT_s_1_3_2((key1[14]), state_1_1_63_32_sva_1_14_1,
          (data_in_rsci_idat_mxwt[14]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_13 <= MUX1HOT_s_1_3_2((key1[13]), state_1_1_63_32_sva_1_13_1,
          (data_in_rsci_idat_mxwt[13]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_12 <= MUX1HOT_s_1_3_2((key1[12]), state_1_1_63_32_sva_1_12_1,
          (data_in_rsci_idat_mxwt[12]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_11 <= MUX1HOT_s_1_3_2((key1[11]), state_1_1_63_32_sva_1_11_1,
          (data_in_rsci_idat_mxwt[11]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_10 <= MUX1HOT_s_1_3_2((key1[10]), state_1_1_63_32_sva_1_10_1,
          (data_in_rsci_idat_mxwt[10]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_9 <= MUX1HOT_s_1_3_2((key1[9]), state_1_1_63_32_sva_1_9_1,
          (data_in_rsci_idat_mxwt[9]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_8 <= MUX1HOT_s_1_3_2((key1[8]), state_1_1_63_32_sva_1_8_1,
          (data_in_rsci_idat_mxwt[8]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_7 <= MUX1HOT_s_1_3_2((key1[7]), state_1_1_63_32_sva_1_7_1,
          (data_in_rsci_idat_mxwt[7]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_6 <= MUX1HOT_s_1_3_2((key1[6]), state_1_1_63_32_sva_1_6_1,
          (data_in_rsci_idat_mxwt[6]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_5 <= MUX1HOT_s_1_3_2((key1[5]), state_1_1_63_32_sva_1_5_1,
          (data_in_rsci_idat_mxwt[5]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_4 <= MUX1HOT_s_1_3_2((key1[4]), state_1_1_63_32_sva_1_4_1,
          (data_in_rsci_idat_mxwt[4]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_3 <= MUX1HOT_s_1_3_2((key1[3]), state_1_1_63_32_sva_1_3_1,
          (data_in_rsci_idat_mxwt[3]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_2 <= MUX1HOT_s_1_3_2((key1[2]), state_1_1_63_32_sva_1_2_1,
          (data_in_rsci_idat_mxwt[2]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_1 <= MUX1HOT_s_1_3_2((key1[1]), state_1_1_63_32_sva_1_1_1,
          (data_in_rsci_idat_mxwt[1]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
      plaintext_63_32_sva_0 <= MUX1HOT_s_1_3_2((key1[0]), state_1_1_63_32_sva_1_0_1,
          (data_in_rsci_idat_mxwt[0]), {(fsm_output[0]) , (fsm_output[1]) , (fsm_output[9])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ADLEN_i_7_0_sva_6_4 <= 3'b000;
      ADLEN_i_7_0_sva_3_0 <= 4'b0000;
    end
    else if ( rst ) begin
      ADLEN_i_7_0_sva_6_4 <= 3'b000;
      ADLEN_i_7_0_sva_3_0 <= 4'b0000;
    end
    else if ( ADLEN_i_and_ssc ) begin
      ADLEN_i_7_0_sva_6_4 <= (z_out_2[6:4]) & (signext_3_1(~ (fsm_output[8]))) &
          (signext_3_1(~ and_740_cse));
      ADLEN_i_7_0_sva_3_0 <= MUX_v_4_2_2(4'b0000, ADLEN_i_ADLEN_i_mux_nl, nor_28_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_1_1_31_0_lpi_4_0 <= 1'b0;
      state_1_1_31_0_lpi_4_1 <= 1'b0;
      state_1_1_31_0_lpi_4_2 <= 1'b0;
      state_1_1_31_0_lpi_4_3 <= 1'b0;
      state_1_1_31_0_lpi_4_4 <= 1'b0;
      state_1_1_31_0_lpi_4_5 <= 1'b0;
      state_1_1_31_0_lpi_4_6 <= 1'b0;
      state_1_1_31_0_lpi_4_7 <= 1'b0;
      state_1_1_31_0_lpi_4_10 <= 1'b0;
      state_1_1_31_0_lpi_4_25 <= 1'b0;
      state_1_1_31_0_lpi_4_26 <= 1'b0;
      state_1_1_31_0_lpi_4_27 <= 1'b0;
      state_1_1_31_0_lpi_4_28 <= 1'b0;
      state_1_1_31_0_lpi_4_29 <= 1'b0;
      state_1_1_31_0_lpi_4_30 <= 1'b0;
      state_1_1_31_0_lpi_4_31 <= 1'b0;
    end
    else if ( rst ) begin
      state_1_1_31_0_lpi_4_0 <= 1'b0;
      state_1_1_31_0_lpi_4_1 <= 1'b0;
      state_1_1_31_0_lpi_4_2 <= 1'b0;
      state_1_1_31_0_lpi_4_3 <= 1'b0;
      state_1_1_31_0_lpi_4_4 <= 1'b0;
      state_1_1_31_0_lpi_4_5 <= 1'b0;
      state_1_1_31_0_lpi_4_6 <= 1'b0;
      state_1_1_31_0_lpi_4_7 <= 1'b0;
      state_1_1_31_0_lpi_4_10 <= 1'b0;
      state_1_1_31_0_lpi_4_25 <= 1'b0;
      state_1_1_31_0_lpi_4_26 <= 1'b0;
      state_1_1_31_0_lpi_4_27 <= 1'b0;
      state_1_1_31_0_lpi_4_28 <= 1'b0;
      state_1_1_31_0_lpi_4_29 <= 1'b0;
      state_1_1_31_0_lpi_4_30 <= 1'b0;
      state_1_1_31_0_lpi_4_31 <= 1'b0;
    end
    else if ( state_and_128_cse ) begin
      state_1_1_31_0_lpi_4_0 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_0_1, state_xor_466_nl,
          state_xor_467_nl, xor_136_nl, state_xor_468_nl, state_3_16_sva_3_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_1 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_1_1, state_xor_470_nl,
          state_xor_471_nl, xor_134_nl, state_xor_472_nl, state_3_17_sva_3_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_2 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_2_1, state_xor_474_nl,
          state_xor_475_nl, xor_132_nl, state_xor_476_nl, state_3_27_sva_3_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_3 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_3_1, state_xor_478_nl,
          state_xor_479_nl, xor_130_nl, state_xor_480_nl, state_3_9_sva_3_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_4 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_4_1, state_xor_482_nl,
          state_xor_483_nl, xor_128_nl, state_xor_484_nl, state_4_60_sva_2_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_5 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_5_1, state_xor_486_nl,
          state_xor_487_nl, xor_126_nl, state_xor_488_nl, state_4_61_sva_2_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_6 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_6_1, state_xor_490_nl,
          state_xor_491_nl, xor_124_nl, state_xor_492_nl, state_4_62_sva_2_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_7 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_7_1, state_xor_494_nl,
          state_xor_495_nl, xor_122_nl, state_xor_496_nl, state_4_63_sva_2_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_10 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_10_1, state_xor_498_nl,
          state_xor_499_nl, xor_116_nl, state_xor_500_nl, state_3_18_sva_3_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_25 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_25_1, state_xor_544_nl,
          state_xor_545_nl, xor_86_nl, state_xor_546_nl, state_3_4_sva_3_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_26 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_26_1, state_xor_548_nl,
          state_xor_549_nl, xor_84_nl, state_xor_550_nl, state_3_5_sva_3_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_27 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_27_1, state_xor_552_nl,
          state_xor_553_nl, xor_82_nl, state_xor_554_nl, state_3_6_sva_3_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_28 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_28_1, state_xor_556_nl,
          state_xor_557_nl, xor_80_nl, state_xor_558_nl, state_3_7_sva_3_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_29 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_29_1, state_xor_560_nl,
          state_xor_561_nl, xor_78_nl, state_xor_562_nl, state_3_8_sva_3_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_30 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_30_1, state_xor_564_nl,
          state_xor_565_nl, xor_76_nl, state_xor_566_nl, state_4_58_sva_2_mx0w5,
          {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse
          , and_94_cse});
      state_1_1_31_0_lpi_4_31 <= MUX1HOT_s_1_6_2(state_1_1_31_0_sva_1_31_1, state_xor_568_nl,
          state_xor_569_nl, xor_5_nl, state_xor_570_nl, state_4_59_sva_2_mx0w5, {(fsm_output[1])
          , (fsm_output[4]) , (fsm_output[11]) , and_885_cse , and_39_cse , and_94_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_1_1_31_0_lpi_4_11 <= 1'b0;
      state_1_1_31_0_lpi_4_12 <= 1'b0;
      state_1_1_31_0_lpi_4_13 <= 1'b0;
      state_1_1_31_0_lpi_4_14 <= 1'b0;
      state_1_1_31_0_lpi_4_15 <= 1'b0;
      state_1_1_31_0_lpi_4_16 <= 1'b0;
      state_1_1_31_0_lpi_4_17 <= 1'b0;
      state_1_1_31_0_lpi_4_18 <= 1'b0;
      state_1_1_31_0_lpi_4_19 <= 1'b0;
      state_1_1_31_0_lpi_4_20 <= 1'b0;
      state_1_1_31_0_lpi_4_21 <= 1'b0;
      state_1_1_31_0_lpi_4_22 <= 1'b0;
      state_1_1_31_0_lpi_4_23 <= 1'b0;
      state_1_1_31_0_lpi_4_24 <= 1'b0;
    end
    else if ( rst ) begin
      state_1_1_31_0_lpi_4_11 <= 1'b0;
      state_1_1_31_0_lpi_4_12 <= 1'b0;
      state_1_1_31_0_lpi_4_13 <= 1'b0;
      state_1_1_31_0_lpi_4_14 <= 1'b0;
      state_1_1_31_0_lpi_4_15 <= 1'b0;
      state_1_1_31_0_lpi_4_16 <= 1'b0;
      state_1_1_31_0_lpi_4_17 <= 1'b0;
      state_1_1_31_0_lpi_4_18 <= 1'b0;
      state_1_1_31_0_lpi_4_19 <= 1'b0;
      state_1_1_31_0_lpi_4_20 <= 1'b0;
      state_1_1_31_0_lpi_4_21 <= 1'b0;
      state_1_1_31_0_lpi_4_22 <= 1'b0;
      state_1_1_31_0_lpi_4_23 <= 1'b0;
      state_1_1_31_0_lpi_4_24 <= 1'b0;
    end
    else if ( state_and_137_cse ) begin
      state_1_1_31_0_lpi_4_11 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_11_1, state_xor_502_nl,
          xor_114_nl, state_xor_503_nl, state_3_19_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_12 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_12_1, state_xor_505_nl,
          xor_112_nl, state_xor_506_nl, state_3_2_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_13 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_13_1, state_xor_508_nl,
          xor_110_nl, state_xor_509_nl, state_3_20_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_14 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_14_1, state_xor_511_nl,
          xor_108_nl, state_xor_512_nl, state_3_21_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_15 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_15_1, state_xor_514_nl,
          xor_106_nl, state_xor_515_nl, state_3_22_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_16 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_16_1, state_xor_517_nl,
          xor_104_nl, state_xor_518_nl, state_3_23_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_17 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_17_1, state_xor_520_nl,
          xor_102_nl, state_xor_521_nl, state_3_24_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_18 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_18_1, state_xor_523_nl,
          xor_100_nl, state_xor_524_nl, state_3_25_sva_3_mx0w4, {(fsm_output[1])
          , and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_19 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_19_1, state_xor_526_nl,
          xor_98_nl, state_xor_527_nl, state_3_26_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_20 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_20_1, state_xor_529_nl,
          xor_96_nl, state_xor_530_nl, state_3_28_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_21 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_21_1, state_xor_532_nl,
          xor_94_nl, state_xor_533_nl, state_3_29_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_22 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_22_1, state_xor_535_nl,
          xor_92_nl, state_xor_536_nl, state_3_3_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_23 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_23_1, state_xor_538_nl,
          xor_90_nl, state_xor_539_nl, state_3_30_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
      state_1_1_31_0_lpi_4_24 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_24_1, state_xor_541_nl,
          xor_88_nl, state_xor_542_nl, state_3_31_sva_3_mx0w4, {(fsm_output[1]) ,
          and_24_cse , and_885_cse , and_39_cse , and_94_cse});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_1_1_31_0_lpi_4_8 <= 1'b0;
      state_1_1_31_0_lpi_4_9 <= 1'b0;
      state_1_1_63_32_lpi_4_0 <= 1'b0;
    end
    else if ( rst ) begin
      state_1_1_31_0_lpi_4_8 <= 1'b0;
      state_1_1_31_0_lpi_4_9 <= 1'b0;
      state_1_1_63_32_lpi_4_0 <= 1'b0;
    end
    else if ( state_and_158_cse ) begin
      state_1_1_31_0_lpi_4_8 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_8_1, state_xor_572_nl,
          state_xor_573_nl, xor_75_nl, state_xor_574_nl, {(fsm_output[1]) , (fsm_output[4])
          , (fsm_output[11]) , and_885_cse , (fsm_output[14])});
      state_1_1_31_0_lpi_4_9 <= MUX1HOT_s_1_5_2(state_1_1_31_0_sva_1_9_1, state_xor_575_nl,
          state_xor_576_nl, xor_77_nl, state_xor_577_nl, {(fsm_output[1]) , (fsm_output[4])
          , (fsm_output[11]) , and_885_cse , (fsm_output[14])});
      state_1_1_63_32_lpi_4_0 <= MUX1HOT_s_1_5_2(state_1_1_63_32_sva_1_0_1, state_xor_578_nl,
          state_xor_579_nl, xor_79_nl, state_xor_580_nl, {(fsm_output[1]) , (fsm_output[4])
          , (fsm_output[11]) , and_885_cse , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_1_1_63_32_lpi_4_1 <= 1'b0;
      state_1_1_63_32_lpi_4_10 <= 1'b0;
      state_1_1_63_32_lpi_4_11 <= 1'b0;
      state_1_1_63_32_lpi_4_12 <= 1'b0;
      state_1_1_63_32_lpi_4_13 <= 1'b0;
      state_1_1_63_32_lpi_4_14 <= 1'b0;
      state_1_1_63_32_lpi_4_15 <= 1'b0;
      state_1_1_63_32_lpi_4_16 <= 1'b0;
      state_1_1_63_32_lpi_4_17 <= 1'b0;
      state_1_1_63_32_lpi_4_18 <= 1'b0;
      state_1_1_63_32_lpi_4_19 <= 1'b0;
      state_1_1_63_32_lpi_4_2 <= 1'b0;
      state_1_1_63_32_lpi_4_20 <= 1'b0;
      state_1_1_63_32_lpi_4_21 <= 1'b0;
      state_1_1_63_32_lpi_4_22 <= 1'b0;
      state_1_1_63_32_lpi_4_23 <= 1'b0;
      state_1_1_63_32_lpi_4_24 <= 1'b0;
      state_1_1_63_32_lpi_4_25 <= 1'b0;
      state_1_1_63_32_lpi_4_26 <= 1'b0;
      state_1_1_63_32_lpi_4_27 <= 1'b0;
      state_1_1_63_32_lpi_4_28 <= 1'b0;
      state_1_1_63_32_lpi_4_29 <= 1'b0;
      state_1_1_63_32_lpi_4_3 <= 1'b0;
      state_1_1_63_32_lpi_4_30 <= 1'b0;
      state_1_1_63_32_lpi_4_31 <= 1'b0;
      state_1_1_63_32_lpi_4_4 <= 1'b0;
      state_1_1_63_32_lpi_4_5 <= 1'b0;
      state_1_1_63_32_lpi_4_6 <= 1'b0;
      state_1_1_63_32_lpi_4_7 <= 1'b0;
      state_1_1_63_32_lpi_4_8 <= 1'b0;
      state_1_1_63_32_lpi_4_9 <= 1'b0;
    end
    else if ( rst ) begin
      state_1_1_63_32_lpi_4_1 <= 1'b0;
      state_1_1_63_32_lpi_4_10 <= 1'b0;
      state_1_1_63_32_lpi_4_11 <= 1'b0;
      state_1_1_63_32_lpi_4_12 <= 1'b0;
      state_1_1_63_32_lpi_4_13 <= 1'b0;
      state_1_1_63_32_lpi_4_14 <= 1'b0;
      state_1_1_63_32_lpi_4_15 <= 1'b0;
      state_1_1_63_32_lpi_4_16 <= 1'b0;
      state_1_1_63_32_lpi_4_17 <= 1'b0;
      state_1_1_63_32_lpi_4_18 <= 1'b0;
      state_1_1_63_32_lpi_4_19 <= 1'b0;
      state_1_1_63_32_lpi_4_2 <= 1'b0;
      state_1_1_63_32_lpi_4_20 <= 1'b0;
      state_1_1_63_32_lpi_4_21 <= 1'b0;
      state_1_1_63_32_lpi_4_22 <= 1'b0;
      state_1_1_63_32_lpi_4_23 <= 1'b0;
      state_1_1_63_32_lpi_4_24 <= 1'b0;
      state_1_1_63_32_lpi_4_25 <= 1'b0;
      state_1_1_63_32_lpi_4_26 <= 1'b0;
      state_1_1_63_32_lpi_4_27 <= 1'b0;
      state_1_1_63_32_lpi_4_28 <= 1'b0;
      state_1_1_63_32_lpi_4_29 <= 1'b0;
      state_1_1_63_32_lpi_4_3 <= 1'b0;
      state_1_1_63_32_lpi_4_30 <= 1'b0;
      state_1_1_63_32_lpi_4_31 <= 1'b0;
      state_1_1_63_32_lpi_4_4 <= 1'b0;
      state_1_1_63_32_lpi_4_5 <= 1'b0;
      state_1_1_63_32_lpi_4_6 <= 1'b0;
      state_1_1_63_32_lpi_4_7 <= 1'b0;
      state_1_1_63_32_lpi_4_8 <= 1'b0;
      state_1_1_63_32_lpi_4_9 <= 1'b0;
    end
    else if ( state_and_161_cse ) begin
      state_1_1_63_32_lpi_4_1 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_1_1, state_xor_581_nl,
          xor_81_nl, state_xor_582_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_10 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_10_1, state_xor_583_nl,
          xor_83_nl, state_xor_584_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_11 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_11_1, state_xor_585_nl,
          xor_85_nl, state_xor_586_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_12 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_12_1, state_xor_587_nl,
          xor_87_nl, state_xor_588_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_13 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_13_1, state_xor_589_nl,
          xor_89_nl, state_xor_590_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_14 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_14_1, state_xor_591_nl,
          xor_91_nl, state_xor_592_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_15 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_15_1, state_xor_593_nl,
          xor_93_nl, state_xor_594_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_16 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_16_1, state_xor_595_nl,
          xor_95_nl, state_xor_596_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_17 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_17_1, state_xor_597_nl,
          xor_97_nl, state_xor_598_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_18 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_18_1, state_xor_599_nl,
          xor_99_nl, state_xor_600_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_19 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_19_1, state_xor_601_nl,
          xor_101_nl, state_xor_602_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_2 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_2_1, state_xor_603_nl,
          xor_103_nl, state_xor_604_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_20 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_20_1, state_xor_605_nl,
          xor_105_nl, state_xor_606_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_21 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_21_1, state_xor_607_nl,
          xor_107_nl, state_xor_608_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_22 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_22_1, state_xor_609_nl,
          xor_109_nl, state_xor_610_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_23 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_23_1, state_xor_611_nl,
          xor_111_nl, state_xor_612_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_24 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_24_1, state_xor_613_nl,
          xor_113_nl, state_xor_614_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_25 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_25_1, state_xor_615_nl,
          xor_115_nl, state_xor_616_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_26 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_26_1, state_xor_617_nl,
          xor_117_nl, state_xor_618_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_27 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_27_1, state_xor_619_nl,
          xor_119_nl, state_xor_620_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_28 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_28_1, state_xor_621_nl,
          xor_121_nl, state_xor_622_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_29 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_29_1, state_xor_623_nl,
          xor_123_nl, state_xor_624_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_3 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_3_1, state_xor_625_nl,
          xor_125_nl, state_xor_626_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_30 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_30_1, state_xor_627_nl,
          xor_127_nl, state_xor_628_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_31 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_31_1, state_xor_629_nl,
          xor_129_nl, state_xor_630_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_4 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_4_1, state_xor_631_nl,
          xor_131_nl, state_xor_632_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_5 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_5_1, state_xor_633_nl,
          xor_133_nl, state_xor_634_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_6 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_6_1, state_xor_635_nl,
          xor_135_nl, state_xor_636_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_7 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_7_1, state_xor_637_nl,
          xor_137_nl, state_xor_638_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_8 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_8_1, state_xor_639_nl,
          xor_120_nl, state_xor_640_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
      state_1_1_63_32_lpi_4_9 <= MUX1HOT_s_1_4_2(state_1_1_63_32_sva_1_9_1, state_xor_641_nl,
          xor_118_nl, state_xor_642_nl, {(fsm_output[1]) , and_24_cse , and_885_cse
          , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_3_0_lpi_3 <= 1'b0;
      state_3_1_lpi_3 <= 1'b0;
      state_3_2_lpi_3 <= 1'b0;
      state_3_3_lpi_3 <= 1'b0;
      state_3_4_lpi_3 <= 1'b0;
      state_3_5_lpi_3 <= 1'b0;
      state_3_6_lpi_3 <= 1'b0;
      state_3_7_lpi_3 <= 1'b0;
      state_3_47_lpi_3 <= 1'b0;
      state_3_48_lpi_3 <= 1'b0;
      state_3_49_lpi_3 <= 1'b0;
      state_3_50_lpi_3 <= 1'b0;
      state_3_51_lpi_3 <= 1'b0;
      state_3_52_lpi_3 <= 1'b0;
      state_3_53_lpi_3 <= 1'b0;
      state_3_54_lpi_3 <= 1'b0;
      state_3_55_lpi_3 <= 1'b0;
      state_3_56_lpi_3 <= 1'b0;
      state_3_57_lpi_3 <= 1'b0;
      state_3_58_lpi_3 <= 1'b0;
      state_3_59_lpi_3 <= 1'b0;
      state_3_60_lpi_3 <= 1'b0;
      state_3_61_lpi_3 <= 1'b0;
    end
    else if ( rst ) begin
      state_3_0_lpi_3 <= 1'b0;
      state_3_1_lpi_3 <= 1'b0;
      state_3_2_lpi_3 <= 1'b0;
      state_3_3_lpi_3 <= 1'b0;
      state_3_4_lpi_3 <= 1'b0;
      state_3_5_lpi_3 <= 1'b0;
      state_3_6_lpi_3 <= 1'b0;
      state_3_7_lpi_3 <= 1'b0;
      state_3_47_lpi_3 <= 1'b0;
      state_3_48_lpi_3 <= 1'b0;
      state_3_49_lpi_3 <= 1'b0;
      state_3_50_lpi_3 <= 1'b0;
      state_3_51_lpi_3 <= 1'b0;
      state_3_52_lpi_3 <= 1'b0;
      state_3_53_lpi_3 <= 1'b0;
      state_3_54_lpi_3 <= 1'b0;
      state_3_55_lpi_3 <= 1'b0;
      state_3_56_lpi_3 <= 1'b0;
      state_3_57_lpi_3 <= 1'b0;
      state_3_58_lpi_3 <= 1'b0;
      state_3_59_lpi_3 <= 1'b0;
      state_3_60_lpi_3 <= 1'b0;
      state_3_61_lpi_3 <= 1'b0;
    end
    else if ( state_and_192_cse ) begin
      state_3_0_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_643_nl, state_xor_644_nl, state_xor_645_nl,
          state_3_0_sva_3_mx0w6, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_1_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_646_nl, state_xor_647_nl, state_xor_648_nl,
          state_3_1_sva_3_mx0w6, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_2_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_649_nl, state_xor_650_nl, state_xor_651_nl,
          state_3_2_sva_3_mx0w4, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_3_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_652_nl, state_xor_653_nl, state_xor_654_nl,
          state_3_3_sva_3_mx0w4, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_4_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_655_nl, state_xor_656_nl, state_xor_657_nl,
          state_3_4_sva_3_mx0w5, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_5_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_658_nl, state_xor_659_nl, state_xor_660_nl,
          state_3_5_sva_3_mx0w5, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_6_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_661_nl, state_xor_662_nl, state_xor_663_nl,
          state_3_6_sva_3_mx0w5, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_7_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_664_nl, state_xor_665_nl, state_xor_666_nl,
          state_3_7_sva_3_mx0w5, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_47_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_769_nl, state_xor_770_nl, state_xor_771_nl,
          state_xor_772_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_48_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_773_nl, state_xor_774_nl, state_xor_775_nl,
          state_xor_776_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_49_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_777_nl, state_xor_778_nl, state_xor_779_nl,
          state_xor_780_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_50_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_781_nl, state_xor_782_nl, state_xor_783_nl,
          state_xor_784_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_51_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_785_nl, state_xor_786_nl, state_xor_787_nl,
          state_xor_788_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_52_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_789_nl, state_xor_790_nl, state_xor_791_nl,
          state_xor_792_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_53_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_793_nl, state_xor_794_nl, state_xor_795_nl,
          state_xor_796_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_54_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_797_nl, state_xor_798_nl, state_xor_799_nl,
          state_xor_800_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_55_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_801_nl, state_xor_802_nl, state_xor_803_nl,
          state_xor_804_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_56_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_805_nl, state_xor_806_nl, state_xor_807_nl,
          state_xor_808_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_57_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_809_nl, state_xor_810_nl, state_xor_811_nl,
          state_xor_812_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_58_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_813_nl, state_xor_814_nl, state_xor_815_nl,
          state_xor_816_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_59_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_817_nl, state_xor_818_nl, state_xor_819_nl,
          state_xor_820_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_60_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_821_nl, state_xor_822_nl, state_xor_823_nl,
          state_xor_824_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
      state_3_61_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_825_nl, state_xor_826_nl, state_xor_827_nl,
          state_xor_828_nl, {(fsm_output[1]) , (fsm_output[4]) , (fsm_output[11])
          , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_4_4_0_lpi_3 <= 1'b0;
    end
    else if ( rst ) begin
      state_4_4_0_lpi_3 <= 1'b0;
    end
    else if ( run_wen & ((fsm_output[1]) | and_24_cse | (fsm_output[8]) | (fsm_output[14]))
        ) begin
      state_4_4_0_lpi_3 <= MUX1HOT_s_1_4_2(state_xor_667_nl, state_xor_668_nl, (~
          state_4_4_0_lpi_3), state_4_0_sva_3, {(fsm_output[1]) , and_24_cse , (fsm_output[8])
          , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_4_4_1_lpi_3 <= 1'b0;
      state_4_4_2_lpi_3 <= 1'b0;
      state_4_4_3_lpi_3 <= 1'b0;
      state_4_4_4_lpi_3 <= 1'b0;
      state_4_4_5_lpi_3 <= 1'b0;
      state_4_4_6_lpi_3 <= 1'b0;
      state_4_4_7_lpi_3 <= 1'b0;
      state_3_15_lpi_3 <= 1'b0;
      state_3_16_lpi_3 <= 1'b0;
      state_3_17_lpi_3 <= 1'b0;
      state_3_18_lpi_3 <= 1'b0;
      state_3_19_lpi_3 <= 1'b0;
      state_3_20_lpi_3 <= 1'b0;
      state_3_21_lpi_3 <= 1'b0;
      state_3_22_lpi_3 <= 1'b0;
      state_3_23_lpi_3 <= 1'b0;
      state_3_24_lpi_3 <= 1'b0;
      state_3_25_lpi_3 <= 1'b0;
      state_3_26_lpi_3 <= 1'b0;
      state_3_27_lpi_3 <= 1'b0;
      state_3_28_lpi_3 <= 1'b0;
      state_3_29_lpi_3 <= 1'b0;
      state_3_30_lpi_3 <= 1'b0;
      state_3_31_lpi_3 <= 1'b0;
      state_3_32_lpi_3 <= 1'b0;
      state_3_33_lpi_3 <= 1'b0;
      state_3_34_lpi_3 <= 1'b0;
      state_3_35_lpi_3 <= 1'b0;
      state_3_36_lpi_3 <= 1'b0;
      state_3_37_lpi_3 <= 1'b0;
      state_3_38_lpi_3 <= 1'b0;
      state_3_39_lpi_3 <= 1'b0;
      state_3_40_lpi_3 <= 1'b0;
      state_3_41_lpi_3 <= 1'b0;
      state_3_42_lpi_3 <= 1'b0;
      state_3_43_lpi_3 <= 1'b0;
      state_3_44_lpi_3 <= 1'b0;
      state_3_45_lpi_3 <= 1'b0;
      state_3_46_lpi_3 <= 1'b0;
      state_3_62_lpi_3 <= 1'b0;
      state_3_63_lpi_3 <= 1'b0;
      state_3_8_lpi_3 <= 1'b0;
      state_3_9_lpi_3 <= 1'b0;
      state_4_4_10_lpi_3 <= 1'b0;
      state_4_4_11_lpi_3 <= 1'b0;
      state_4_4_12_lpi_3 <= 1'b0;
      state_4_4_13_lpi_3 <= 1'b0;
      state_4_4_14_lpi_3 <= 1'b0;
      state_4_4_15_lpi_3 <= 1'b0;
      state_4_4_16_lpi_3 <= 1'b0;
      state_4_4_17_lpi_3 <= 1'b0;
      state_4_4_18_lpi_3 <= 1'b0;
      state_4_4_19_lpi_3 <= 1'b0;
      state_4_4_20_lpi_3 <= 1'b0;
      state_4_4_21_lpi_3 <= 1'b0;
      state_4_4_22_lpi_3 <= 1'b0;
      state_4_4_25_lpi_3 <= 1'b0;
      state_4_4_26_lpi_3 <= 1'b0;
      state_4_4_27_lpi_3 <= 1'b0;
      state_4_4_28_lpi_3 <= 1'b0;
      state_4_4_29_lpi_3 <= 1'b0;
      state_4_4_30_lpi_3 <= 1'b0;
      state_4_4_31_lpi_3 <= 1'b0;
      state_4_4_32_lpi_3 <= 1'b0;
      state_4_4_33_lpi_3 <= 1'b0;
      state_4_4_34_lpi_3 <= 1'b0;
      state_4_4_35_lpi_3 <= 1'b0;
      state_4_4_36_lpi_3 <= 1'b0;
      state_4_4_37_lpi_3 <= 1'b0;
      state_4_4_38_lpi_3 <= 1'b0;
      state_4_4_39_lpi_3 <= 1'b0;
      state_4_4_40_lpi_3 <= 1'b0;
      state_4_4_41_lpi_3 <= 1'b0;
      state_4_4_42_lpi_3 <= 1'b0;
      state_4_4_43_lpi_3 <= 1'b0;
      state_4_4_44_lpi_3 <= 1'b0;
      state_4_4_45_lpi_3 <= 1'b0;
      state_4_4_46_lpi_3 <= 1'b0;
      state_4_4_47_lpi_3 <= 1'b0;
      state_4_4_48_lpi_3 <= 1'b0;
      state_4_4_49_lpi_3 <= 1'b0;
      state_4_4_50_lpi_3 <= 1'b0;
      state_4_4_51_lpi_3 <= 1'b0;
      state_4_4_52_lpi_3 <= 1'b0;
      state_4_4_53_lpi_3 <= 1'b0;
      state_4_4_54_lpi_3 <= 1'b0;
      state_4_4_55_lpi_3 <= 1'b0;
      state_4_4_56_lpi_3 <= 1'b0;
      state_4_4_57_lpi_3 <= 1'b0;
      state_4_4_58_lpi_3 <= 1'b0;
      state_4_4_59_lpi_3 <= 1'b0;
      state_4_4_60_lpi_3 <= 1'b0;
      state_4_4_61_lpi_3 <= 1'b0;
      state_4_4_62_lpi_3 <= 1'b0;
      state_4_4_63_lpi_3 <= 1'b0;
      state_4_4_8_lpi_3 <= 1'b0;
      state_4_4_9_lpi_3 <= 1'b0;
    end
    else if ( rst ) begin
      state_4_4_1_lpi_3 <= 1'b0;
      state_4_4_2_lpi_3 <= 1'b0;
      state_4_4_3_lpi_3 <= 1'b0;
      state_4_4_4_lpi_3 <= 1'b0;
      state_4_4_5_lpi_3 <= 1'b0;
      state_4_4_6_lpi_3 <= 1'b0;
      state_4_4_7_lpi_3 <= 1'b0;
      state_3_15_lpi_3 <= 1'b0;
      state_3_16_lpi_3 <= 1'b0;
      state_3_17_lpi_3 <= 1'b0;
      state_3_18_lpi_3 <= 1'b0;
      state_3_19_lpi_3 <= 1'b0;
      state_3_20_lpi_3 <= 1'b0;
      state_3_21_lpi_3 <= 1'b0;
      state_3_22_lpi_3 <= 1'b0;
      state_3_23_lpi_3 <= 1'b0;
      state_3_24_lpi_3 <= 1'b0;
      state_3_25_lpi_3 <= 1'b0;
      state_3_26_lpi_3 <= 1'b0;
      state_3_27_lpi_3 <= 1'b0;
      state_3_28_lpi_3 <= 1'b0;
      state_3_29_lpi_3 <= 1'b0;
      state_3_30_lpi_3 <= 1'b0;
      state_3_31_lpi_3 <= 1'b0;
      state_3_32_lpi_3 <= 1'b0;
      state_3_33_lpi_3 <= 1'b0;
      state_3_34_lpi_3 <= 1'b0;
      state_3_35_lpi_3 <= 1'b0;
      state_3_36_lpi_3 <= 1'b0;
      state_3_37_lpi_3 <= 1'b0;
      state_3_38_lpi_3 <= 1'b0;
      state_3_39_lpi_3 <= 1'b0;
      state_3_40_lpi_3 <= 1'b0;
      state_3_41_lpi_3 <= 1'b0;
      state_3_42_lpi_3 <= 1'b0;
      state_3_43_lpi_3 <= 1'b0;
      state_3_44_lpi_3 <= 1'b0;
      state_3_45_lpi_3 <= 1'b0;
      state_3_46_lpi_3 <= 1'b0;
      state_3_62_lpi_3 <= 1'b0;
      state_3_63_lpi_3 <= 1'b0;
      state_3_8_lpi_3 <= 1'b0;
      state_3_9_lpi_3 <= 1'b0;
      state_4_4_10_lpi_3 <= 1'b0;
      state_4_4_11_lpi_3 <= 1'b0;
      state_4_4_12_lpi_3 <= 1'b0;
      state_4_4_13_lpi_3 <= 1'b0;
      state_4_4_14_lpi_3 <= 1'b0;
      state_4_4_15_lpi_3 <= 1'b0;
      state_4_4_16_lpi_3 <= 1'b0;
      state_4_4_17_lpi_3 <= 1'b0;
      state_4_4_18_lpi_3 <= 1'b0;
      state_4_4_19_lpi_3 <= 1'b0;
      state_4_4_20_lpi_3 <= 1'b0;
      state_4_4_21_lpi_3 <= 1'b0;
      state_4_4_22_lpi_3 <= 1'b0;
      state_4_4_25_lpi_3 <= 1'b0;
      state_4_4_26_lpi_3 <= 1'b0;
      state_4_4_27_lpi_3 <= 1'b0;
      state_4_4_28_lpi_3 <= 1'b0;
      state_4_4_29_lpi_3 <= 1'b0;
      state_4_4_30_lpi_3 <= 1'b0;
      state_4_4_31_lpi_3 <= 1'b0;
      state_4_4_32_lpi_3 <= 1'b0;
      state_4_4_33_lpi_3 <= 1'b0;
      state_4_4_34_lpi_3 <= 1'b0;
      state_4_4_35_lpi_3 <= 1'b0;
      state_4_4_36_lpi_3 <= 1'b0;
      state_4_4_37_lpi_3 <= 1'b0;
      state_4_4_38_lpi_3 <= 1'b0;
      state_4_4_39_lpi_3 <= 1'b0;
      state_4_4_40_lpi_3 <= 1'b0;
      state_4_4_41_lpi_3 <= 1'b0;
      state_4_4_42_lpi_3 <= 1'b0;
      state_4_4_43_lpi_3 <= 1'b0;
      state_4_4_44_lpi_3 <= 1'b0;
      state_4_4_45_lpi_3 <= 1'b0;
      state_4_4_46_lpi_3 <= 1'b0;
      state_4_4_47_lpi_3 <= 1'b0;
      state_4_4_48_lpi_3 <= 1'b0;
      state_4_4_49_lpi_3 <= 1'b0;
      state_4_4_50_lpi_3 <= 1'b0;
      state_4_4_51_lpi_3 <= 1'b0;
      state_4_4_52_lpi_3 <= 1'b0;
      state_4_4_53_lpi_3 <= 1'b0;
      state_4_4_54_lpi_3 <= 1'b0;
      state_4_4_55_lpi_3 <= 1'b0;
      state_4_4_56_lpi_3 <= 1'b0;
      state_4_4_57_lpi_3 <= 1'b0;
      state_4_4_58_lpi_3 <= 1'b0;
      state_4_4_59_lpi_3 <= 1'b0;
      state_4_4_60_lpi_3 <= 1'b0;
      state_4_4_61_lpi_3 <= 1'b0;
      state_4_4_62_lpi_3 <= 1'b0;
      state_4_4_63_lpi_3 <= 1'b0;
      state_4_4_8_lpi_3 <= 1'b0;
      state_4_4_9_lpi_3 <= 1'b0;
    end
    else if ( state_and_201_cse ) begin
      state_4_4_1_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_670_nl, state_xor_671_nl, state_4_1_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_2_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_673_nl, state_xor_674_nl, state_4_2_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_3_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_675_nl, state_xor_676_nl, state_4_3_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_4_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_677_nl, state_xor_678_nl, state_4_4_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_5_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_679_nl, state_xor_680_nl, state_4_5_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_6_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_681_nl, state_xor_682_nl, state_4_6_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_7_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_683_nl, state_xor_684_nl, state_4_7_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_15_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_690_nl, state_xor_691_nl, state_3_15_sva_3_mx0w6,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_16_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_692_nl, state_xor_693_nl, state_3_16_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_17_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_694_nl, state_xor_695_nl, state_3_17_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_18_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_696_nl, state_xor_697_nl, state_3_18_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_19_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_698_nl, state_xor_699_nl, state_3_19_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_20_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_700_nl, state_xor_701_nl, state_3_20_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_21_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_702_nl, state_xor_703_nl, state_3_21_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_22_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_704_nl, state_xor_705_nl, state_3_22_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_23_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_706_nl, state_xor_707_nl, state_3_23_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_24_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_708_nl, state_xor_709_nl, state_3_24_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_25_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_710_nl, state_xor_711_nl, state_3_25_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_26_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_712_nl, state_xor_713_nl, state_3_26_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_27_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_714_nl, state_xor_715_nl, state_3_27_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_28_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_716_nl, state_xor_717_nl, state_3_28_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_29_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_718_nl, state_xor_719_nl, state_3_29_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_30_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_720_nl, state_xor_721_nl, state_3_30_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_31_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_722_nl, state_xor_723_nl, state_3_31_sva_3_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_32_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_724_nl, state_xor_725_nl, state_xor_726_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_33_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_727_nl, state_xor_728_nl, state_xor_729_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_34_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_730_nl, state_xor_731_nl, state_xor_732_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_35_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_733_nl, state_xor_734_nl, state_xor_735_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_36_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_736_nl, state_xor_737_nl, state_xor_738_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_37_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_739_nl, state_xor_740_nl, state_xor_741_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_38_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_742_nl, state_xor_743_nl, state_xor_744_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_39_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_745_nl, state_xor_746_nl, state_xor_747_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_40_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_748_nl, state_xor_749_nl, state_xor_750_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_41_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_751_nl, state_xor_752_nl, state_xor_753_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_42_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_754_nl, state_xor_755_nl, state_xor_756_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_43_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_757_nl, state_xor_758_nl, state_xor_759_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_44_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_760_nl, state_xor_761_nl, state_xor_762_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_45_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_763_nl, state_xor_764_nl, state_xor_765_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_46_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_766_nl, state_xor_767_nl, state_xor_768_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_62_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_829_nl, state_xor_830_nl, state_xor_831_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_63_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_832_nl, state_xor_833_nl, state_xor_834_nl,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_8_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_835_nl, state_xor_836_nl, state_3_8_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_3_9_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_837_nl, state_xor_838_nl, state_3_9_sva_3_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_10_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_839_nl, state_xor_840_nl, state_4_10_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_11_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_842_nl, state_xor_843_nl, state_4_11_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_12_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_845_nl, state_xor_846_nl, state_4_12_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_13_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_848_nl, state_xor_849_nl, state_4_13_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_14_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_851_nl, state_xor_852_nl, state_4_14_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_15_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_854_nl, state_xor_855_nl, state_4_15_sva_3,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_16_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_857_nl, state_xor_858_nl, state_4_16_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_17_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_859_nl, state_xor_860_nl, state_4_17_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_18_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_861_nl, state_xor_862_nl, state_4_18_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_19_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_863_nl, state_xor_864_nl, state_4_19_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_20_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_865_nl, state_xor_866_nl, state_4_20_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_21_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_867_nl, state_xor_868_nl, state_4_21_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_22_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_869_nl, state_xor_870_nl, state_4_22_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_25_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_873_nl, state_xor_874_nl, state_4_25_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_26_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_875_nl, state_xor_876_nl, state_4_26_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_27_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_877_nl, state_xor_878_nl, state_4_27_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_28_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_879_nl, state_xor_880_nl, state_4_28_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_29_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_881_nl, state_xor_882_nl, state_4_29_sva_2_mx0w4,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_30_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_883_nl, state_xor_884_nl, state_4_30_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_31_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_885_nl, state_xor_886_nl, state_4_31_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_32_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_887_nl, state_xor_888_nl, state_4_32_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_33_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_889_nl, state_xor_890_nl, state_4_33_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_34_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_891_nl, state_xor_892_nl, state_4_34_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_35_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_893_nl, state_xor_894_nl, state_4_35_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_36_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_895_nl, state_xor_896_nl, state_4_36_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_37_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_897_nl, state_xor_898_nl, state_4_37_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_38_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_899_nl, state_xor_900_nl, state_4_38_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_39_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_901_nl, state_xor_902_nl, state_4_39_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_40_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_903_nl, state_xor_904_nl, state_4_40_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_41_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_905_nl, state_xor_906_nl, state_4_41_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_42_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_907_nl, state_xor_908_nl, state_4_42_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_43_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_909_nl, state_xor_910_nl, state_4_43_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_44_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_911_nl, state_xor_912_nl, state_4_44_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_45_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_913_nl, state_xor_914_nl, state_4_45_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_46_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_915_nl, state_xor_916_nl, state_4_46_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_47_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_917_nl, state_xor_918_nl, state_4_47_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_48_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_919_nl, state_xor_920_nl, state_4_48_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_49_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_921_nl, state_xor_922_nl, state_4_49_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_50_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_923_nl, state_xor_924_nl, state_4_50_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_51_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_925_nl, state_xor_926_nl, state_4_51_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_52_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_927_nl, state_xor_928_nl, state_4_52_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_53_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_929_nl, state_xor_930_nl, state_4_53_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_54_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_931_nl, state_xor_932_nl, state_4_54_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_55_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_933_nl, state_xor_934_nl, state_4_55_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_56_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_935_nl, state_xor_936_nl, state_4_56_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_57_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_937_nl, state_xor_938_nl, state_4_57_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_58_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_939_nl, state_xor_940_nl, state_4_58_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_59_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_941_nl, state_xor_942_nl, state_4_59_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_60_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_943_nl, state_xor_944_nl, state_4_60_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_61_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_945_nl, state_xor_946_nl, state_4_61_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_62_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_947_nl, state_xor_948_nl, state_4_62_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_63_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_949_nl, state_xor_950_nl, state_4_63_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_8_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_951_nl, state_xor_952_nl, state_4_8_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
      state_4_4_9_lpi_3 <= MUX1HOT_s_1_3_2(state_xor_953_nl, state_xor_954_nl, state_4_9_sva_2_mx0w5,
          {(fsm_output[1]) , and_24_cse , (fsm_output[14])});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_3_10_lpi_3 <= 1'b0;
      state_3_11_lpi_3 <= 1'b0;
      state_3_12_lpi_3 <= 1'b0;
      state_3_13_lpi_3 <= 1'b0;
      state_3_14_lpi_3 <= 1'b0;
      state_4_4_23_lpi_3 <= 1'b0;
      state_4_4_24_lpi_3 <= 1'b0;
    end
    else if ( rst ) begin
      state_3_10_lpi_3 <= 1'b0;
      state_3_11_lpi_3 <= 1'b0;
      state_3_12_lpi_3 <= 1'b0;
      state_3_13_lpi_3 <= 1'b0;
      state_3_14_lpi_3 <= 1'b0;
      state_4_4_23_lpi_3 <= 1'b0;
      state_4_4_24_lpi_3 <= 1'b0;
    end
    else if ( state_and_208_cse ) begin
      state_3_10_lpi_3 <= MUX_s_1_2_2(state_xor_685_nl, state_3_10_sva_2_mx0w6, or_tmp_1693);
      state_3_11_lpi_3 <= MUX_s_1_2_2(state_xor_686_nl, state_3_11_sva_2_mx0w6, or_tmp_1693);
      state_3_12_lpi_3 <= MUX_s_1_2_2(state_xor_687_nl, state_3_12_sva_2_mx0w6, or_tmp_1693);
      state_3_13_lpi_3 <= MUX_s_1_2_2(state_xor_688_nl, state_3_13_sva_2_mx0w6, or_tmp_1693);
      state_3_14_lpi_3 <= MUX_s_1_2_2(state_xor_689_nl, state_3_14_sva_2_mx0w6, or_tmp_1693);
      state_4_4_23_lpi_3 <= MUX_s_1_2_2(state_xor_871_nl, state_4_4_23_sva_1_mx0w4,
          or_tmp_1693);
      state_4_4_24_lpi_3 <= MUX_s_1_2_2(state_xor_872_nl, state_4_4_24_sva_1_mx0w4,
          or_tmp_1693);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_2_0_1_lpi_6 <= 1'b0;
      state_2_1_1_lpi_6 <= 1'b0;
      state_2_2_1_lpi_6 <= 1'b0;
      state_2_3_1_lpi_6 <= 1'b0;
      state_2_4_1_lpi_6 <= 1'b0;
      state_2_5_1_lpi_6 <= 1'b0;
      state_2_6_1_lpi_6 <= 1'b0;
      state_2_7_1_lpi_6 <= 1'b0;
    end
    else if ( rst ) begin
      state_2_0_1_lpi_6 <= 1'b0;
      state_2_1_1_lpi_6 <= 1'b0;
      state_2_2_1_lpi_6 <= 1'b0;
      state_2_3_1_lpi_6 <= 1'b0;
      state_2_4_1_lpi_6 <= 1'b0;
      state_2_5_1_lpi_6 <= 1'b0;
      state_2_6_1_lpi_6 <= 1'b0;
      state_2_7_1_lpi_6 <= 1'b0;
    end
    else if ( state_and_320_cse ) begin
      state_2_0_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_0_1_sva_4, state_xnor_176_nl,
          state_4_0_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_1_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_1_1_sva_4, state_xnor_177_nl,
          state_4_1_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_2_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_2_1_sva_4, state_xnor_178_nl,
          state_4_10_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_3_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_3_1_sva_4, state_xnor_179_nl,
          state_4_11_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_4_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_4_1_sva_4, state_xnor_180_nl,
          state_4_12_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_5_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_5_1_sva_4, state_xnor_181_nl,
          state_4_13_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_6_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_6_1_sva_4, state_xnor_182_nl,
          state_4_14_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
      state_2_7_1_lpi_6 <= MUX1HOT_s_1_3_2(state_2_7_1_sva_4, state_xnor_183_nl,
          state_4_15_sva_3, {(fsm_output[4]) , (fsm_output[11]) , (fsm_output[14])});
    end
  end
  assign PLEN_xor_62_nl = plaintext_31_0_sva_0 ^ state_0_0_lpi_6;
  assign xor_403_nl = xor_cse_7 ^ xor_cse_10 ^ xor_cse_11 ^ xor_cse_12 ^ state_1_1_31_0_lpi_4_8
      ^ state_1_1_63_32_lpi_4_16 ^ (key1[0]);
  assign xor_262_nl = state_2_0_1_lpi_4 ^ (key2[0]);
  assign PLEN_xor_60_nl = plaintext_31_0_sva_1 ^ state_0_1_lpi_6;
  assign xor_418_nl = xor_cse_21 ^ xor_cse_24 ^ xor_cse_25 ^ xor_cse_26 ^ state_1_1_31_0_lpi_4_9
      ^ state_1_1_63_32_lpi_4_17 ^ (key1[1]);
  assign xor_260_nl = state_2_1_1_lpi_4 ^ (key2[1]);
  assign PLEN_xor_58_nl = plaintext_31_0_sva_2 ^ state_0_2_lpi_6;
  assign xor_432_nl = xor_cse_34 ^ xor_cse_37 ^ xor_cse_38 ^ xor_cse_39 ^ Encrypt_Top_sbox_2_and_750
      ^ state_1_1_63_32_lpi_4_0 ^ (key1[2]);
  assign xor_258_nl = state_1_1_31_0_lpi_4_12 ^ (key2[2]);
  assign xor_321_nl = state_2_14_1_lpi_4 ^ (key4[2]);
  assign PLEN_xor_56_nl = plaintext_31_0_sva_3 ^ state_0_3_lpi_6;
  assign xor_447_nl = xor_cse_48 ^ xor_cse_51 ^ xor_cse_52 ^ xor_cse_53 ^ state_1_1_63_32_lpi_4_1
      ^ state_1_1_63_32_lpi_4_19 ^ (key1[3]);
  assign xor_256_nl = state_1_1_31_0_lpi_4_22 ^ (key2[3]);
  assign xor_319_nl = state_2_25_1_lpi_4 ^ (key4[3]);
  assign PLEN_xor_54_nl = plaintext_31_0_sva_4 ^ state_0_32_lpi_6;
  assign xor_462_nl = xor_cse_62 ^ xor_cse_65 ^ xor_cse_66 ^ xor_cse_67 ^ state_1_1_63_32_lpi_4_10
      ^ state_1_1_63_32_lpi_4_2 ^ (key1[4]);
  assign xor_254_nl = state_1_1_31_0_lpi_4_25 ^ (key2[4]);
  assign xor_317_nl = state_2_28_1_lpi_4 ^ (key4[4]);
  assign PLEN_xor_52_nl = plaintext_31_0_sva_5 ^ state_0_33_lpi_6;
  assign xor_477_nl = xor_cse_76 ^ xor_cse_79 ^ xor_cse_80 ^ xor_cse_81 ^ state_1_1_63_32_lpi_4_11
      ^ state_1_1_63_32_lpi_4_20 ^ (key1[5]);
  assign xor_252_nl = state_1_1_31_0_lpi_4_26 ^ (key2[5]);
  assign xor_315_nl = state_2_29_1_lpi_4 ^ (key4[5]);
  assign PLEN_xor_50_nl = plaintext_31_0_sva_6 ^ state_0_34_lpi_6;
  assign xor_492_nl = xor_cse_90 ^ xor_cse_94 ^ xor_cse_95 ^ Encrypt_Top_sbox_2_and_636
      ^ Encrypt_Top_sbox_2_and_638 ^ state_1_1_63_32_lpi_4_21 ^ (key1[6]);
  assign xor_250_nl = state_1_1_31_0_lpi_4_27 ^ (key2[6]);
  assign xor_313_nl = state_2_30_1_lpi_4 ^ (key4[6]);
  assign PLEN_xor_48_nl = plaintext_31_0_sva_7 ^ state_0_35_lpi_6;
  assign xor_506_nl = xor_cse_104 ^ xor_cse_106 ^ xor_cse_107 ^ xor_cse_108 ^ state_1_1_63_32_lpi_4_13
      ^ state_1_1_63_32_lpi_4_22 ^ (key1[7]);
  assign xor_248_nl = state_1_1_31_0_lpi_4_28 ^ (key2[7]);
  assign xor_311_nl = state_2_31_1_lpi_4 ^ (key4[7]);
  assign PLEN_xor_46_nl = plaintext_31_0_sva_8 ^ state_0_36_lpi_6;
  assign xor_520_nl = xor_cse_117 ^ xor_cse_119 ^ xor_cse_120 ^ xor_cse_121 ^ state_1_1_63_32_lpi_4_14
      ^ state_1_1_63_32_lpi_4_23 ^ (key1[8]);
  assign xor_246_nl = state_1_1_31_0_lpi_4_29 ^ (key2[8]);
  assign PLEN_xor_44_nl = plaintext_31_0_sva_9 ^ state_0_37_lpi_6;
  assign xor_533_nl = xor_cse_129 ^ xor_cse_132 ^ xor_cse_37 ^ xor_cse_133 ^ state_1_1_63_32_lpi_4_15
      ^ state_1_1_63_32_lpi_4_24 ^ (key1[9]);
  assign xor_244_nl = state_1_1_31_0_lpi_4_3 ^ (key2[9]);
  assign PLEN_xor_42_nl = plaintext_31_0_sva_10 ^ state_0_10_lpi_6;
  assign xor_546_nl = xor_cse_141 ^ xor_cse_143 ^ xor_cse_145 ^ state_1_1_63_32_lpi_4_25
      ^ (key1[10]);
  assign xor_242_nl = state_2_2_1_lpi_4 ^ (key2[10]);
  assign xor_305_nl = state_2_2_1_lpi_6 ^ (key4[10]);
  assign PLEN_xor_40_nl = plaintext_31_0_sva_11 ^ state_0_11_lpi_6;
  assign xor_558_nl = xor_cse_153 ^ xor_cse_65 ^ xor_cse_22 ^ xor_cse_156 ^ Encrypt_Top_sbox_2_and_598
      ^ state_1_1_63_32_lpi_4_26 ^ (key1[11]);
  assign xor_240_nl = state_2_3_1_lpi_4 ^ (key2[11]);
  assign xor_303_nl = state_2_3_1_lpi_6 ^ (key4[11]);
  assign PLEN_xor_38_nl = plaintext_31_0_sva_12 ^ state_0_12_lpi_6;
  assign xor_568_nl = xor_cse_34 ^ xor_cse_163 ^ xor_cse_79 ^ state_1_1_63_32_lpi_4_27
      ^ Encrypt_Top_sbox_2_and_532 ^ state_1_1_63_32_lpi_4_5 ^ (key1[12]);
  assign xor_238_nl = state_2_4_1_lpi_4 ^ (key2[12]);
  assign xor_301_nl = state_2_4_1_lpi_6 ^ (key4[12]);
  assign PLEN_xor_36_nl = plaintext_31_0_sva_13 ^ state_0_13_lpi_6;
  assign xor_579_nl = xor_cse_172 ^ xor_cse_174 ^ xor_cse_49 ^ xor_cse_175 ^ Encrypt_Top_sbox_2_and_662
      ^ state_1_1_63_32_lpi_4_19 ^ (key1[13]);
  assign xor_236_nl = state_2_5_1_lpi_4 ^ (key2[13]);
  assign xor_299_nl = state_2_5_1_lpi_6 ^ (key4[13]);
  assign PLEN_xor_34_nl = plaintext_31_0_sva_14 ^ state_0_14_lpi_6;
  assign xor_591_nl = xor_cse_183 ^ xor_cse_185 ^ xor_cse_63 ^ xor_cse_186 ^ Encrypt_Top_sbox_2_and_654
      ^ state_1_1_63_32_lpi_4_2 ^ (key1[14]);
  assign xor_234_nl = state_2_6_1_lpi_4 ^ (key2[14]);
  assign xor_297_nl = state_2_6_1_lpi_6 ^ (key4[14]);
  assign PLEN_xor_nl = plaintext_31_0_sva_15 ^ state_0_15_lpi_6;
  assign xor_604_nl = xor_cse_194 ^ xor_cse_195 ^ xor_cse_77 ^ state_1_1_63_32_lpi_4_3
      ^ (key1[15]);
  assign xor_232_nl = state_2_7_1_lpi_4 ^ (key2[15]);
  assign xor_295_nl = state_2_7_1_lpi_6 ^ (key4[15]);
  assign PLEN_xor_33_nl = plaintext_31_0_sva_16 ^ state_0_16_lpi_6;
  assign xor_615_nl = xor_cse_205 ^ (key1[16]) ^ xor_cse_132 ^ xor_cse_94 ^ xor_cse_209;
  assign xor_230_nl = state_1_1_31_0_lpi_4_0 ^ (key2[16]);
  assign xor_293_nl = state_2_10_1_lpi_4 ^ (key4[16]);
  assign PLEN_xor_35_nl = plaintext_31_0_sva_17 ^ state_0_17_lpi_6;
  assign xor_626_nl = xor_cse_141 ^ xor_cse_217 ^ xor_cse_10 ^ xor_cse_218 ^ Encrypt_Top_sbox_2_and_628
      ^ Encrypt_Top_sbox_2_and_630 ^ state_1_1_63_32_lpi_4_22 ^ (key1[17]);
  assign xor_228_nl = state_1_1_31_0_lpi_4_1 ^ (key2[17]);
  assign xor_291_nl = state_2_11_1_lpi_4 ^ (key4[17]);
  assign PLEN_xor_37_nl = plaintext_31_0_sva_18 ^ state_0_18_lpi_6;
  assign xor_637_nl = xor_cse_153 ^ xor_cse_226 ^ (key1[18]) ^ xor_cse_228 ^ xor_cse_229;
  assign xor_226_nl = state_1_1_31_0_lpi_4_10 ^ (key2[18]);
  assign xor_289_nl = state_2_12_1_lpi_4 ^ (key4[18]);
  assign PLEN_xor_39_nl = plaintext_31_0_sva_19 ^ state_0_19_lpi_6;
  assign xor_649_nl = xor_cse_235 ^ xor_cse_238 ^ xor_cse_239 ^ state_1_1_63_32_lpi_4_5
      ^ (key1[19]);
  assign xor_224_nl = state_1_1_31_0_lpi_4_11 ^ (key2[19]);
  assign xor_287_nl = state_2_13_1_lpi_4 ^ (key4[19]);
  assign PLEN_xor_41_nl = plaintext_31_0_sva_20 ^ state_0_20_lpi_6;
  assign xor_660_nl = xor_cse_246 ^ xor_cse_248 ^ xor_cse_51 ^ xor_cse_249 ^ Encrypt_Top_sbox_2_and_606
      ^ state_1_1_63_32_lpi_4_25 ^ state_1_1_63_32_lpi_4_6 ^ (key1[20]);
  assign xor_222_nl = state_1_1_31_0_lpi_4_13 ^ (key2[20]);
  assign xor_285_nl = state_2_15_1_lpi_4 ^ (key4[20]);
  assign PLEN_xor_43_nl = plaintext_31_0_sva_21 ^ state_0_21_lpi_6;
  assign xor_672_nl = xor_cse_256 ^ xor_cse_257 ^ xor_cse_260 ^ state_1_1_63_32_lpi_4_7
      ^ (key1[21]);
  assign xor_220_nl = state_1_1_31_0_lpi_4_14 ^ (key2[21]);
  assign xor_283_nl = state_2_16_1_lpi_4 ^ (key4[21]);
  assign PLEN_xor_45_nl = plaintext_31_0_sva_22 ^ state_0_22_lpi_6;
  assign xor_683_nl = xor_cse_267 ^ xor_cse_196 ^ xor_cse_197 ^ xor_cse_270 ^ state_1_1_63_32_lpi_4_27
      ^ (key1[22]);
  assign xor_218_nl = state_1_1_31_0_lpi_4_15 ^ (key2[22]);
  assign xor_281_nl = state_2_17_1_lpi_4 ^ (key4[22]);
  assign PLEN_xor_47_nl = plaintext_31_0_sva_23 ^ state_0_23_lpi_6;
  assign xor_692_nl = xor_cse_277 ^ xor_cse_172 ^ (key1[23]) ^ xor_cse_206 ^ xor_cse_207;
  assign xor_216_nl = state_1_1_31_0_lpi_4_16 ^ (key2[23]);
  assign xor_279_nl = state_2_18_1_lpi_4 ^ (key4[23]);
  assign PLEN_xor_49_nl = plaintext_31_0_sva_24 ^ state_0_24_lpi_6;
  assign xor_701_nl = xor_cse_183 ^ xor_cse_285 ^ (key1[24]) ^ xor_cse_217 ^ xor_cse_218;
  assign xor_214_nl = state_1_1_31_0_lpi_4_17 ^ (key2[24]);
  assign xor_277_nl = state_2_19_1_lpi_4 ^ (key4[24]);
  assign PLEN_xor_51_nl = plaintext_31_0_sva_25 ^ state_0_25_lpi_6;
  assign xor_711_nl = xor_cse_293 ^ xor_cse_228 ^ xor_cse_229 ^ state_1_1_63_32_lpi_4_3
      ^ (key1[25]);
  assign xor_212_nl = state_1_1_31_0_lpi_4_18 ^ (key2[25]);
  assign xor_275_nl = state_2_20_1_lpi_4 ^ (key4[25]);
  assign PLEN_xor_53_nl = plaintext_31_0_sva_26 ^ state_0_26_lpi_6;
  assign xor_721_nl = xor_cse_302 ^ xor_cse_238 ^ xor_cse_239 ^ state_1_1_63_32_lpi_4_30
      ^ (key1[26]);
  assign xor_210_nl = state_1_1_31_0_lpi_4_19 ^ (key2[26]);
  assign xor_316_nl = state_1_1_31_0_lpi_4_30 ^ (key3[26]);
  assign xor_273_nl = state_2_21_1_lpi_4 ^ (key4[26]);
  assign PLEN_xor_55_nl = plaintext_31_0_sva_27 ^ state_0_27_lpi_6;
  assign xor_731_nl = xor_cse_311 ^ xor_cse_248 ^ xor_cse_249 ^ state_1_1_63_32_lpi_4_31
      ^ (key1[27]);
  assign xor_208_nl = state_1_1_31_0_lpi_4_2 ^ (key2[27]);
  assign xor_318_nl = state_1_1_31_0_lpi_4_31 ^ (key3[27]);
  assign xor_271_nl = state_2_22_1_lpi_4 ^ (key4[27]);
  assign PLEN_xor_57_nl = plaintext_31_0_sva_28 ^ state_0_28_lpi_6;
  assign xor_741_nl = xor_cse_320 ^ xor_cse_258 ^ xor_cse_260 ^ state_1_1_63_32_lpi_4_4
      ^ (key1[28]);
  assign xor_206_nl = state_1_1_31_0_lpi_4_20 ^ (key2[28]);
  assign xor_320_nl = state_1_1_31_0_lpi_4_4 ^ (key3[28]);
  assign xor_269_nl = state_2_23_1_lpi_4 ^ (key4[28]);
  assign PLEN_xor_59_nl = plaintext_31_0_sva_29 ^ state_0_29_lpi_6;
  assign xor_751_nl = xor_cse_329 ^ xor_cse_270 ^ xor_cse_331 ^ state_1_1_63_32_lpi_4_5
      ^ (key1[29]);
  assign xor_204_nl = state_1_1_31_0_lpi_4_21 ^ (key2[29]);
  assign xor_322_nl = state_1_1_31_0_lpi_4_5 ^ (key3[29]);
  assign xor_267_nl = state_2_24_1_lpi_4 ^ (key4[29]);
  assign PLEN_xor_61_nl = plaintext_31_0_sva_30 ^ state_0_30_lpi_6;
  assign xor_760_nl = xor_cse_277 ^ xor_cse_174 ^ xor_cse_231 ^ xor_cse_339 ^ Encrypt_Top_sbox_2_and_526
      ^ state_1_1_63_32_lpi_4_6 ^ (key1[30]);
  assign xor_202_nl = state_1_1_31_0_lpi_4_23 ^ (key2[30]);
  assign xor_324_nl = state_1_1_31_0_lpi_4_6 ^ (key3[30]);
  assign xor_265_nl = state_2_26_1_lpi_4 ^ (key4[30]);
  assign PLEN_xor_63_nl = plaintext_31_0_sva_31 ^ state_0_31_lpi_6;
  assign xor_769_nl = xor_cse_285 ^ xor_cse_185 ^ xor_cse_242 ^ xor_cse_347 ^ Encrypt_Top_sbox_2_and_518
      ^ state_1_1_63_32_lpi_4_7 ^ (key1[31]);
  assign xor_9_nl = state_1_1_31_0_lpi_4_24 ^ (key2[31]);
  assign xor_326_nl = state_1_1_31_0_lpi_4_7 ^ (key3[31]);
  assign xor_11_nl = state_2_27_1_lpi_4 ^ (key4[31]);
  assign state_xor_338_nl = xor_cse_1731 ^ xor_cse_1732 ^ xor_cse_1733;
  assign state_xor_340_nl = xor_cse_1739 ^ xor_cse_1097 ^ xor_cse_1740;
  assign state_xor_342_nl = xor_cse_1087 ^ xor_cse_1746 ^ xor_cse_1747;
  assign state_xor_344_nl = xor_cse_1078 ^ xor_cse_1753 ^ xor_cse_1754;
  assign state_xor_346_nl = xor_cse_1752 ^ xor_cse_1758 ^ xor_cse_1759;
  assign state_xor_348_nl = xor_cse_1745 ^ xor_cse_1763 ^ xor_cse_1764;
  assign state_xor_350_nl = xor_cse_1738 ^ xor_cse_1768 ^ xor_cse_1769;
  assign state_xor_352_nl = xor_cse_1773 ^ xor_cse_1732 ^ xor_cse_1774;
  assign state_xor_354_nl = xor_cse_1097 ^ xor_cse_1778 ^ xor_cse_1779;
  assign state_xor_356_nl = xor_cse_1087 ^ xor_cse_1783 ^ xor_cse_1784;
  assign state_xor_358_nl = xor_cse_1078 ^ xor_cse_1787 ^ xor_cse_1788;
  assign state_xor_360_nl = xor_cse_1792 ^ xor_cse_1758 ^ xor_cse_1793;
  assign state_xor_362_nl = xor_cse_1789 ^ xor_cse_1763 ^ xor_cse_1795;
  assign state_xor_364_nl = xor_cse_1785 ^ xor_cse_1768 ^ xor_cse_1797;
  assign state_xor_366_nl = xor_cse_1773 ^ xor_cse_1781 ^ xor_cse_1799;
  assign state_xor_368_nl = xor_cse_1776 ^ xor_cse_1778 ^ xor_cse_1801;
  assign state_xor_370_nl = xor_cse_1771 ^ xor_cse_1783 ^ xor_cse_1803;
  assign state_xor_372_nl = xor_cse_403 ^ xor_cse_1766 ^ xor_cse_1787 ^ Encrypt_Top_sbox_and_2_cse_46_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_53_sva_1 ^ state_4_3_31_0_sva_23;
  assign state_xor_374_nl = xor_cse_1761 ^ xor_cse_387 ^ xor_cse_1792 ^ Encrypt_Top_sbox_and_2_cse_45_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_52_sva_1 ^ state_4_3_31_0_sva_22;
  assign state_xor_376_nl = xor_cse_1756 ^ xor_cse_375 ^ xor_cse_1789 ^ Encrypt_Top_sbox_and_2_cse_44_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_51_sva_1 ^ state_4_3_31_0_sva_21;
  assign state_xor_378_nl = xor_cse_1749 ^ xor_cse_362 ^ xor_cse_1785 ^ Encrypt_Top_sbox_and_2_cse_43_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_50_sva_1 ^ state_4_3_31_0_sva_20;
  assign state_xor_380_nl = xor_cse_1742 ^ xor_cse_350 ^ xor_cse_1781 ^ Encrypt_Top_sbox_and_2_cse_42_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_49_sva_1 ^ state_4_3_31_0_sva_19;
  assign state_xor_382_nl = xor_cse_1736 ^ xor_cse_951 ^ xor_cse_1776 ^ Encrypt_Top_sbox_and_2_cse_41_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_48_sva_1 ^ state_4_3_31_0_sva_18;
  assign state_xor_384_nl = xor_cse_1731 ^ xor_cse_1771 ^ xor_cse_1790 ^ Encrypt_Top_sbox_and_2_cse_40_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_47_sva_1 ^ Encrypt_Top_sbox_and_2_cse_17_sva_1;
  assign state_xor_386_nl = xor_cse_1739 ^ xor_cse_926 ^ xor_cse_1766 ^ Encrypt_Top_sbox_and_2_cse_39_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_46_sva_1 ^ state_4_3_31_0_sva_16;
  assign state_xor_388_nl = xor_cse_1761 ^ xor_cse_912 ^ xor_cse_1746 ^ Encrypt_Top_sbox_and_2_cse_38_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_45_sva_1 ^ state_4_3_31_0_sva_15;
  assign state_xor_390_nl = xor_cse_1756 ^ xor_cse_900 ^ xor_cse_1753 ^ Encrypt_Top_sbox_and_2_cse_37_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_44_sva_1 ^ state_4_3_31_0_sva_14;
  assign state_xor_392_nl = xor_cse_1749 ^ xor_cse_890 ^ xor_cse_1760 ^ Encrypt_Top_sbox_and_2_cse_36_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_43_sva_1 ^ state_4_3_31_0_sva_13;
  assign state_xor_394_nl = xor_cse_1742 ^ xor_cse_880 ^ xor_cse_1765 ^ Encrypt_Top_sbox_and_2_cse_35_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_42_sva_1 ^ state_4_3_31_0_sva_12;
  assign state_xor_396_nl = xor_cse_1736 ^ xor_cse_868 ^ xor_cse_1770 ^ Encrypt_Top_sbox_and_2_cse_34_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_41_sva_1 ^ state_4_3_31_0_sva_11;
  assign state_xor_398_nl = xor_cse_1731 ^ xor_cse_861 ^ xor_cse_1775 ^ Encrypt_Top_sbox_and_2_cse_33_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_40_sva_1 ^ state_4_3_31_0_sva_10;
  assign state_xor_400_nl = xor_cse_1739 ^ xor_cse_1780 ^ xor_cse_1750 ^ Encrypt_Top_sbox_and_2_cse_32_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_39_sva_1 ^ Encrypt_Top_sbox_and_2_cse_9_sva_1;
  assign state_xor_402_nl = xor_cse_1835 ^ xor_cse_1838 ^ xor_cse_1172 ^ xor_cse_1842;
  assign state_xor_404_nl = xor_cse_1855 ^ xor_cse_1162 ^ xor_cse_1400 ^ xor_cse_1859
      ^ xor_cse_1864 ^ state_4_3_31_0_sva_8;
  assign state_xor_406_nl = xor_cse_444 ^ xor_cse_1874 ^ xor_cse_1877 ^ xor_cse_1880;
  assign state_xor_408_nl = xor_cse_430 ^ xor_cse_1892 ^ xor_cse_1895 ^ xor_cse_1898;
  assign state_xor_410_nl = xor_cse_417 ^ xor_cse_1907 ^ xor_cse_1886 ^ xor_cse_1910;
  assign state_xor_412_nl = xor_cse_405 ^ xor_cse_1913 ^ xor_cse_1868 ^ xor_cse_1919;
  assign state_xor_414_nl = xor_cse_389 ^ xor_cse_1901 ^ xor_cse_1845 ^ xor_cse_1925;
  assign state_xor_416_nl = xor_cse_1931 ^ xor_cse_377 ^ xor_cse_1172 ^ xor_cse_1883
      ^ xor_cse_1842;
  assign state_xor_418_nl = xor_cse_1941 ^ xor_cse_364 ^ xor_cse_1162 ^ xor_cse_1865
      ^ xor_cse_1945;
  assign state_xor_420_nl = xor_cse_1951 ^ xor_cse_352 ^ xor_cse_444 ^ xor_cse_1849
      ^ xor_cse_1874;
  assign state_xor_422_nl = xor_cse_430 ^ xor_cse_1892 ^ xor_cse_1838 ^ xor_cse_1960;
  assign state_xor_424_nl = xor_cse_417 ^ xor_cse_1907 ^ xor_cse_1966 ^ xor_cse_1969;
  assign state_xor_426_nl = xor_cse_405 ^ xor_cse_1913 ^ xor_cse_1973 ^ xor_cse_1880;
  assign state_xor_428_nl = xor_cse_389 ^ xor_cse_1901 ^ xor_cse_1979 ^ xor_cse_1898;
  assign state_xor_430_nl = xor_cse_377 ^ xor_cse_1883 ^ xor_cse_1910 ^ xor_cse_1985;
  assign state_xor_432_nl = xor_cse_364 ^ xor_cse_1865 ^ xor_cse_1919 ^ xor_cse_1991;
  assign state_xor_434_nl = xor_cse_352 ^ xor_cse_1849 ^ xor_cse_1925 ^ xor_cse_1998;
  assign state_xor_436_nl = xor_cse_1838 ^ xor_cse_1931 ^ xor_cse_948 ^ xor_cse_2005;
  assign state_xor_438_nl = xor_cse_1941 ^ xor_cse_2013 ^ xor_cse_1969;
  assign state_xor_440_nl = xor_cse_1951 ^ xor_cse_924 ^ xor_cse_1375 ^ xor_cse_2021
      ^ xor_cse_2024 ^ state_4_3_63_32_sva_12;
  assign state_xor_442_nl = xor_cse_1960 ^ xor_cse_910 ^ xor_cse_1528 ^ xor_cse_2029
      ^ xor_cse_2032 ^ state_4_3_63_32_sva_11;
  assign state_xor_444_nl = xor_cse_1910 ^ xor_cse_1966 ^ xor_cse_2036;
  assign state_xor_446_nl = xor_cse_1919 ^ xor_cse_1973 ^ xor_cse_888 ^ xor_cse_2044;
  assign state_xor_448_nl = xor_cse_1925 ^ xor_cse_1979 ^ xor_cse_878 ^ xor_cse_2053;
  assign state_xor_450_nl = xor_cse_1931 ^ xor_cse_1985 ^ xor_cse_2047;
  assign state_xor_452_nl = xor_cse_1941 ^ xor_cse_1991 ^ xor_2162_cse;
  assign state_xor_454_nl = xor_cse_1951 ^ xor_cse_1998 ^ xor_cse_2033;
  assign state_xor_456_nl = xor_cse_1960 ^ xor_cse_2025 ^ xor_2168_cse;
  assign state_xor_458_nl = xor_cse_1966 ^ xor_cse_2013 ^ xor_2172_cse;
  assign state_xor_460_nl = xor_cse_1973 ^ xor_cse_2008 ^ xor_cse_924 ^ xor_cse_2069;
  assign state_xor_462_nl = xor_cse_1979 ^ xor_cse_2001 ^ xor_cse_910 ^ xor_cse_2065;
  assign state_xor_464_nl = xor_cse_2036 ^ xor_cse_1985 ^ xor_2184_cse;
  assign state_xor_401_nl = xor_cse_390 ^ xor_cse_1746 ^ xor_cse_1743 ^ state_4_3_31_0_sva_31
      ^ Encrypt_Top_sbox_and_2_cse_38_sva_1 ^ Encrypt_Top_sbox_and_2_cse_8_sva_1;
  assign state_xor_399_nl = xor_cse_1735 ^ xor_cse_379 ^ xor_cse_1753 ^ state_4_3_31_0_sva_30
      ^ Encrypt_Top_sbox_and_2_cse_37_sva_1 ^ Encrypt_Top_sbox_and_2_cse_7_sva_1;
  assign state_xor_397_nl = xor_cse_1734 ^ xor_cse_366 ^ xor_cse_1760 ^ state_4_3_31_0_sva_29
      ^ Encrypt_Top_sbox_and_2_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_6_sva_1;
  assign state_xor_395_nl = xor_cse_1741 ^ xor_cse_354 ^ xor_cse_1765 ^ state_4_3_31_0_sva_28
      ^ Encrypt_Top_sbox_and_2_cse_35_sva_1 ^ Encrypt_Top_sbox_and_2_cse_5_sva_1;
  assign state_xor_393_nl = xor_cse_1748 ^ xor_cse_1031 ^ xor_cse_1770 ^ state_4_3_31_0_sva_27
      ^ Encrypt_Top_sbox_and_2_cse_34_sva_1 ^ Encrypt_Top_sbox_and_2_cse_4_sva_1;
  assign state_xor_391_nl = xor_cse_1755 ^ xor_cse_448 ^ xor_cse_1775 ^ state_4_3_31_0_sva_26
      ^ Encrypt_Top_sbox_and_2_cse_33_sva_1 ^ Encrypt_Top_sbox_and_2_cse_3_sva_1;
  assign state_xor_389_nl = xor_cse_1752 ^ xor_cse_428 ^ xor_cse_1780 ^ state_4_3_31_0_sva_25
      ^ Encrypt_Top_sbox_and_2_cse_32_sva_1 ^ Encrypt_Top_sbox_and_2_cse_2_sva_1;
  assign state_xor_387_nl = xor_cse_1745 ^ xor_cse_390 ^ xor_cse_415 ^ state_4_3_31_0_sva_24
      ^ state_4_3_31_0_sva_31 ^ Encrypt_Top_sbox_and_2_cse_1_sva_1;
  assign state_xor_385_nl = xor_cse_1738 ^ xor_cse_379 ^ xor_cse_403 ^ state_4_3_31_0_sva_23
      ^ state_4_3_31_0_sva_30 ^ Encrypt_Top_sbox_and_2_cse_0_sva_1;
  assign state_xor_383_nl = xor_cse_366 ^ xor_cse_387 ^ xor_cse_1732 ^ state_4_3_31_0_sva_22
      ^ state_4_3_31_0_sva_29 ^ Encrypt_Top_sbox_and_2_cse_63_sva_1;
  assign state_xor_381_nl = xor_cse_1097 ^ xor_cse_354 ^ xor_cse_375 ^ state_4_3_31_0_sva_21
      ^ state_4_3_31_0_sva_28 ^ state_4_3_63_32_sva_30;
  assign state_xor_379_nl = xor_cse_1087 ^ xor_cse_362 ^ xor_cse_1031 ^ state_4_3_31_0_sva_20
      ^ state_4_3_31_0_sva_27 ^ state_4_3_63_32_sva_29;
  assign state_xor_377_nl = xor_cse_1078 ^ xor_cse_350 ^ xor_cse_448 ^ state_4_3_31_0_sva_19
      ^ state_4_3_31_0_sva_26 ^ state_4_3_63_32_sva_28;
  assign state_xor_375_nl = xor_cse_428 ^ xor_cse_951 ^ xor_cse_1758 ^ state_4_3_31_0_sva_18
      ^ state_4_3_31_0_sva_25 ^ Encrypt_Top_sbox_and_2_cse_59_sva_1;
  assign state_xor_373_nl = xor_cse_415 ^ xor_cse_1790 ^ xor_cse_1763 ^ Encrypt_Top_sbox_and_2_cse_17_sva_1
      ^ state_4_3_31_0_sva_24 ^ Encrypt_Top_sbox_and_2_cse_58_sva_1;
  assign state_xor_371_nl = xor_cse_926 ^ xor_cse_1768 ^ xor_cse_1804;
  assign state_xor_369_nl = xor_cse_1773 ^ xor_cse_912 ^ xor_cse_1802;
  assign state_xor_367_nl = xor_cse_900 ^ xor_cse_1778 ^ xor_cse_1800;
  assign state_xor_365_nl = xor_cse_890 ^ xor_cse_1783 ^ xor_cse_1798;
  assign state_xor_363_nl = xor_cse_880 ^ xor_cse_1787 ^ xor_cse_1796;
  assign state_xor_361_nl = xor_cse_868 ^ xor_cse_1792 ^ xor_cse_1794;
  assign state_xor_359_nl = xor_cse_861 ^ xor_cse_1789 ^ xor_cse_1790 ^ state_4_3_31_0_sva_10
      ^ Encrypt_Top_sbox_and_2_cse_17_sva_1 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1;
  assign state_xor_357_nl = xor_cse_1785 ^ xor_cse_1750 ^ xor_cse_1786;
  assign state_xor_355_nl = xor_cse_1781 ^ xor_cse_1743 ^ xor_cse_1782;
  assign state_xor_353_nl = xor_cse_1735 ^ xor_cse_1776 ^ xor_cse_1777;
  assign state_xor_351_nl = xor_cse_1734 ^ xor_cse_1771 ^ xor_cse_1772;
  assign state_xor_349_nl = xor_cse_1741 ^ xor_cse_1766 ^ xor_cse_1767;
  assign state_xor_347_nl = xor_cse_1748 ^ xor_cse_1761 ^ xor_cse_1762;
  assign state_xor_345_nl = xor_cse_1755 ^ xor_cse_1756 ^ xor_cse_1757;
  assign state_xor_343_nl = xor_cse_1749 ^ xor_cse_1750 ^ xor_cse_1751;
  assign state_xor_341_nl = xor_cse_1742 ^ xor_cse_1743 ^ xor_cse_1744;
  assign state_xor_339_nl = xor_cse_1735 ^ xor_cse_1736 ^ xor_cse_1737;
  assign state_xor_465_nl = xor_cse_1988 ^ xor_cse_1991 ^ xor_2186_cse;
  assign state_xor_463_nl = xor_cse_1982 ^ xor_cse_1998 ^ xor_2182_cse;
  assign state_xor_461_nl = xor_cse_1976 ^ xor_cse_2047 ^ xor_2168_cse;
  assign state_xor_459_nl = xor_cse_1970 ^ xor_cse_2013 ^ xor_2162_cse;
  assign state_xor_457_nl = xor_cse_1963 ^ xor_cse_2033 ^ xor_cse_924 ^ xor_cse_2069;
  assign state_xor_455_nl = xor_cse_1955 ^ xor_cse_2025 ^ xor_cse_910 ^ xor_cse_2065;
  assign state_xor_453_nl = xor_cse_1946 ^ xor_cse_2036 ^ xor_2172_cse;
  assign state_xor_451_nl = xor_cse_1936 ^ xor_cse_2008 ^ xor_2186_cse;
  assign state_xor_449_nl = xor_cse_1928 ^ xor_cse_2001 ^ xor_2182_cse;
  assign state_xor_447_nl = xor_cse_1922 ^ xor_cse_2047 ^ xor_2184_cse;
  assign state_xor_445_nl = xor_cse_1916 ^ xor_cse_1988 ^ xor_cse_859 ^ xor_cse_2040;
  assign state_xor_443_nl = xor_cse_1904 ^ xor_cse_1982 ^ xor_cse_2033;
  assign state_xor_441_nl = xor_cse_1889 ^ xor_cse_1976 ^ xor_cse_2025;
  assign state_xor_439_nl = xor_cse_1871 ^ xor_cse_1970 ^ xor_cse_446 ^ xor_cse_2017;
  assign state_xor_437_nl = xor_cse_1963 ^ xor_cse_2008 ^ xor_cse_933 ^ xor_cse_1852;
  assign state_xor_435_nl = xor_cse_1835 ^ xor_cse_1955 ^ xor_cse_2001;
  assign state_xor_433_nl = xor_cse_1855 ^ xor_cse_1946 ^ xor_cse_401 ^ xor_cse_1995;
  assign state_xor_431_nl = xor_cse_1877 ^ xor_cse_1936 ^ xor_cse_1988;
  assign state_xor_429_nl = xor_cse_1895 ^ xor_cse_1928 ^ xor_cse_1982;
  assign state_xor_427_nl = xor_cse_1886 ^ xor_cse_1922 ^ xor_cse_1976;
  assign state_xor_425_nl = xor_cse_1868 ^ xor_cse_1916 ^ xor_cse_1970;
  assign state_xor_423_nl = xor_cse_1845 ^ xor_cse_1904 ^ xor_cse_1963;
  assign state_xor_421_nl = xor_cse_1889 ^ xor_cse_1955 ^ xor_cse_1172 ^ xor_cse_1842;
  assign state_xor_419_nl = xor_cse_1871 ^ xor_cse_1946 ^ xor_cse_1162 ^ xor_cse_1945;
  assign state_xor_417_nl = xor_cse_1936 ^ xor_cse_444 ^ xor_cse_933 ^ xor_cse_1874
      ^ xor_cse_1852;
  assign state_xor_415_nl = xor_cse_430 ^ xor_cse_1892 ^ xor_cse_1835 ^ xor_cse_1928;
  assign state_xor_413_nl = xor_cse_417 ^ xor_cse_1907 ^ xor_cse_1855 ^ xor_cse_1922;
  assign state_xor_411_nl = xor_cse_405 ^ xor_cse_1913 ^ xor_cse_1877 ^ xor_cse_1916;
  assign state_xor_409_nl = xor_cse_389 ^ xor_cse_1901 ^ xor_cse_1895 ^ xor_cse_1904;
  assign state_xor_407_nl = xor_cse_377 ^ xor_cse_1883 ^ xor_cse_1886 ^ xor_cse_1889;
  assign state_xor_405_nl = xor_cse_364 ^ xor_cse_1865 ^ xor_cse_1868 ^ xor_cse_1871;
  assign state_xor_403_nl = xor_cse_1845 ^ xor_cse_352 ^ xor_cse_933 ^ xor_cse_1849
      ^ xor_cse_1852;
  assign state_xor_nl = xor_cse_349 ^ xor_cse_351 ^ xor_cse_354 ^ plaintext_31_0_sva_0
      ^ Encrypt_Top_sbox_and_1_cse_28_sva_1 ^ state_2_28_1_lpi_4 ^ state_0_28_lpi_6;
  assign state_xor_1_nl = xor_cse_56 ^ xor_cse_356 ^ xor_cse_358 ^ xor_cse_359;
  assign state_xor_2_nl = xor_cse_56 ^ xor_cse_60 ^ xor_cse_356 ^ xor_cse_358;
  assign state_xor_3_nl = xor_cse_56 ^ xor_cse_360 ^ xor_cse_356 ^ xor_cse_358;
  assign mux1h_nl = MUX1HOT_s_1_6_2(state_xor_nl, state_0_0_sva_2_mx0w1, state_xor_1_nl,
      state_xor_2_nl, data_out_rsci_idat_0, state_xor_3_nl, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_4_nl = xor_cse_361 ^ xor_cse_363 ^ xor_cse_366 ^ plaintext_31_0_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_29_sva_1 ^ state_2_29_1_lpi_4 ^ state_0_29_lpi_6;
  assign state_xor_5_nl = xor_cse_368 ^ xor_cse_370 ^ xor_cse_70 ^ Encrypt_Top_sbox_1_and_1_cse_1_sva_1
      ^ state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ state_0_1_lpi_6;
  assign state_xor_6_nl = xor_cse_70 ^ xor_cse_71 ^ xor_cse_368 ^ xor_cse_370;
  assign state_xor_7_nl = xor_cse_70 ^ xor_cse_373 ^ xor_cse_368 ^ xor_cse_370;
  assign mux1h_1_nl = MUX1HOT_s_1_6_2(state_xor_4_nl, state_0_1_sva_2_mx0w1, state_xor_5_nl,
      state_xor_6_nl, data_out_rsci_idat_1, state_xor_7_nl, {(fsm_output[1]) , (fsm_output[3])
      , (fsm_output[4]) , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_8_nl = xor_cse_374 ^ xor_cse_376 ^ xor_cse_379 ^ plaintext_31_0_sva_2
      ^ Encrypt_Top_sbox_and_1_cse_30_sva_1 ^ state_2_30_1_lpi_4 ^ state_0_30_lpi_6;
  assign state_xor_9_nl = xor_cse_84 ^ xor_cse_381 ^ xor_cse_382 ^ xor_cse_383;
  assign state_xor_10_nl = xor_cse_84 ^ xor_cse_88 ^ xor_cse_381 ^ xor_cse_383;
  assign state_xor_11_nl = xor_cse_84 ^ xor_cse_381 ^ xor_cse_383 ^ xor_cse_385;
  assign mux1h_2_nl = MUX1HOT_s_1_6_2(state_xor_8_nl, state_0_2_sva_2_mx0w1, state_xor_9_nl,
      state_xor_10_nl, data_out_rsci_idat_2, state_xor_11_nl, {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_12_nl = xor_cse_386 ^ xor_cse_389 ^ xor_cse_390 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_3
      ^ Encrypt_Top_sbox_and_1_cse_3_sva_1 ^ Encrypt_Top_sbox_and_2_cse_3_sva_1 ^
      plaintext_31_0_sva_3 ^ Encrypt_Top_sbox_and_1_cse_31_sva_1 ^ state_2_31_1_lpi_4
      ^ state_0_31_lpi_6;
  assign state_xor_13_nl = xor_cse_393 ^ xor_cse_395 ^ xor_cse_102 ^ Encrypt_Top_sbox_1_and_1_cse_3_sva_1
      ^ state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3])
      ^ state_0_3_lpi_6;
  assign state_xor_14_nl = xor_cse_102 ^ xor_cse_103 ^ xor_cse_393 ^ xor_cse_395;
  assign state_xor_15_nl = xor_cse_393 ^ xor_cse_395 ^ xor_cse_102 ^ Encrypt_Top_sbox_3_and_1_cse_3_sva_1
      ^ state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ state_0_3_lpi_6;
  assign mux1h_3_nl = MUX1HOT_s_1_6_2(state_xor_12_nl, state_0_3_sva_2_mx0w1, state_xor_13_nl,
      state_xor_14_nl, data_out_rsci_idat_3, state_xor_15_nl, {(fsm_output[1]) ,
      (fsm_output[3]) , (fsm_output[4]) , (fsm_output[11]) , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_16_nl = xor_cse_400 ^ xor_cse_402 ^ xor_cse_405 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_4
      ^ Encrypt_Top_sbox_and_1_cse_4_sva_1 ^ Encrypt_Top_sbox_and_2_cse_4_sva_1 ^
      plaintext_31_0_sva_4;
  assign state_xor_17_nl = xor_cse_407 ^ Encrypt_Top_sbox_1_and_1_cse_32_sva_1 ^
      xor_cse_4 ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1 ^ state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4])
      ^ state_0_4_lpi_6;
  assign state_xor_19_nl = xor_cse_407 ^ Encrypt_Top_sbox_3_and_1_cse_32_sva_1 ^
      xor_cse_412 ^ Encrypt_Top_sbox_3_and_1_cse_4_sva_1 ^ state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4])
      ^ state_0_4_lpi_6;
  assign mux1h_4_nl = MUX1HOT_s_1_7_2(state_xor_16_nl, state_0_4_sva_2_mx0w1, state_xor_17_nl,
      state_0_4_sva_4_mx0w4, ciphertext_32_sva_mx0w2, data_out_rsci_idat_4, state_xor_19_nl,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_20_nl = xor_cse_414 ^ xor_cse_416 ^ xor_cse_419 ^ plaintext_31_0_sva_5
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_1 ^ Encrypt_Top_sbox_and_1_cse_33_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_33_sva_1;
  assign state_xor_21_nl = xor_cse_421 ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1 ^
      xor_cse_18 ^ Encrypt_Top_sbox_1_and_1_cse_5_sva_1 ^ state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5])
      ^ state_0_5_lpi_6;
  assign state_xor_23_nl = Encrypt_Top_sbox_3_and_1_cse_33_sva_1 ^ xor_cse_425 ^
      xor_cse_426 ^ xor_cse_421;
  assign mux1h_5_nl = MUX1HOT_s_1_7_2(state_xor_20_nl, state_0_5_sva_2_mx0w1, state_xor_21_nl,
      state_0_5_sva_4_mx0w4, ciphertext_33_sva_mx0w2, data_out_rsci_idat_5, state_xor_23_nl,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_24_nl = xor_cse_427 ^ xor_cse_430 ^ xor_cse_431 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_6
      ^ Encrypt_Top_sbox_and_1_cse_6_sva_1 ^ Encrypt_Top_sbox_and_2_cse_6_sva_1 ^
      plaintext_31_0_sva_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_2 ^ Encrypt_Top_sbox_and_1_cse_34_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_34_sva_1;
  assign state_xor_25_nl = xor_cse_325 ^ xor_cse_136 ^ xor_cse_30 ^ xor_cse_434 ^
      xor_cse_435 ^ xor_cse_436;
  assign state_xor_27_nl = xor_cse_438 ^ xor_cse_325 ^ xor_cse_136 ^ xor_cse_441
      ^ Encrypt_Top_sbox_1_and_cse_25_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_25_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1;
  assign mux1h_6_nl = MUX1HOT_s_1_7_2(state_xor_24_nl, state_0_6_sva_2_mx0w1, state_xor_25_nl,
      state_0_6_sva_4_mx0w4, ciphertext_34_sva_mx0w2, data_out_rsci_idat_6, state_xor_27_nl,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_28_nl = xor_cse_443 ^ xor_cse_445 ^ xor_cse_448 ^ plaintext_31_0_sva_7
      ^ Encrypt_Top_sbox_and_1_cse_26_sva_1 ^ state_2_26_1_lpi_4 ^ state_0_26_lpi_6;
  assign state_xor_29_nl = xor_cse_450 ^ xor_cse_148 ^ xor_cse_46 ^ xor_cse_452 ^
      xor_cse_453;
  assign state_xor_31_nl = xor_cse_148 ^ xor_cse_456 ^ xor_cse_450 ^ xor_cse_457;
  assign mux1h_7_nl = MUX1HOT_s_1_7_2(state_xor_28_nl, state_0_7_sva_2_mx0w1, state_xor_29_nl,
      state_0_7_sva_4_mx0w4, ciphertext_35_sva_mx0w2, data_out_rsci_idat_7, state_xor_31_nl,
      {(fsm_output[1]) , (fsm_output[3]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[13]) , (fsm_output[14])});
  assign state_xnor_nl = ~(xor_cse_459 ^ xor_cse_461 ^ xor_cse_463);
  assign state_xnor_1_nl = ~(xor_cse_465 ^ xor_cse_466 ^ xor_cse_467);
  assign xor_53_nl = state_2_10_1_lpi_4 ^ (key4[10]);
  assign state_xnor_2_nl = ~(xor_cse_472 ^ xor_cse_463 ^ xor_cse_475);
  assign state_xnor_3_nl = ~(xor_cse_466 ^ xor_cse_477 ^ Encrypt_Top_sbox_1_and_786
      ^ state_4_4_17_lpi_3 ^ state_2_17_1_lpi_4 ^ state_1_1_31_0_lpi_4_17);
  assign xor_51_nl = state_2_11_1_lpi_4 ^ (key4[11]);
  assign state_xnor_4_nl = ~(xor_cse_483 ^ xor_cse_475 ^ xor_cse_487 ^ state_4_3_31_0_sva_13
      ^ state_2_13_1_lpi_4 ^ plaintext_31_0_sva_13);
  assign state_xnor_5_nl = ~(xor_cse_477 ^ xor_cse_488 ^ Encrypt_Top_sbox_1_and_788
      ^ state_4_4_18_lpi_3 ^ state_2_18_1_lpi_4 ^ state_1_1_31_0_lpi_4_18);
  assign xor_49_nl = state_2_12_1_lpi_4 ^ (key4[12]);
  assign state_xnor_6_nl = ~(xor_cse_487 ^ state_4_3_31_0_sva_13 ^ state_2_13_1_lpi_4
      ^ plaintext_31_0_sva_13 ^ xor_cse_494 ^ state_4_3_31_0_sva_14 ^ state_2_14_1_lpi_4
      ^ plaintext_31_0_sva_14 ^ xor_cse_495 ^ state_4_3_31_0_sva_19 ^ state_2_19_1_lpi_4
      ^ plaintext_31_0_sva_19);
  assign state_xnor_7_nl = ~(xor_cse_488 ^ xor_cse_496 ^ Encrypt_Top_sbox_1_and_790
      ^ state_4_4_19_lpi_3 ^ state_2_19_1_lpi_4 ^ state_1_1_31_0_lpi_4_19);
  assign xor_47_nl = state_2_13_1_lpi_4 ^ (key4[13]);
  assign state_xnor_8_nl = ~(xor_cse_494 ^ state_4_3_31_0_sva_14 ^ state_2_14_1_lpi_4
      ^ plaintext_31_0_sva_14 ^ xor_cse_502 ^ state_4_3_31_0_sva_15 ^ state_2_15_1_lpi_4
      ^ plaintext_31_0_sva_15 ^ xor_cse_503 ^ state_4_3_31_0_sva_20 ^ state_2_20_1_lpi_4
      ^ plaintext_31_0_sva_20);
  assign state_xnor_9_nl = ~(xor_cse_504 ^ xor_cse_496 ^ xor_cse_505);
  assign xor_45_nl = state_2_14_1_lpi_4 ^ (key4[14]);
  assign state_xnor_10_nl = ~(xor_cse_459 ^ xor_cse_509 ^ xor_cse_511 ^ state_4_3_31_0_sva_21
      ^ state_2_21_1_lpi_4 ^ plaintext_31_0_sva_21);
  assign state_xnor_11_nl = ~(xor_cse_504 ^ xor_cse_467 ^ xor_cse_513);
  assign xor_43_nl = state_2_15_1_lpi_4 ^ (key4[15]);
  assign state_xnor_12_nl = ~(xor_cse_472 ^ xor_cse_459 ^ xor_cse_519 ^ state_4_3_31_0_sva_22
      ^ state_2_22_1_lpi_4 ^ plaintext_31_0_sva_22);
  assign state_xnor_13_nl = ~(Encrypt_Top_sbox_1_and_784 ^ state_4_4_16_lpi_3 ^ state_2_16_1_lpi_4
      ^ state_1_1_31_0_lpi_4_16 ^ Encrypt_Top_sbox_1_and_786 ^ state_4_4_17_lpi_3
      ^ state_2_17_1_lpi_4 ^ state_1_1_31_0_lpi_4_17 ^ Encrypt_Top_sbox_1_and_796
      ^ state_4_4_22_lpi_3 ^ state_2_22_1_lpi_4 ^ state_1_1_31_0_lpi_4_22);
  assign xor_41_nl = state_2_16_1_lpi_4 ^ (key4[16]);
  assign state_xnor_14_nl = ~(xor_cse_472 ^ xor_cse_483 ^ xor_cse_525 ^ state_4_3_31_0_sva_23
      ^ state_2_23_1_lpi_4 ^ plaintext_31_0_sva_23);
  assign state_xnor_15_nl = ~(Encrypt_Top_sbox_1_and_786 ^ state_4_4_17_lpi_3 ^ state_2_17_1_lpi_4
      ^ state_1_1_31_0_lpi_4_17 ^ Encrypt_Top_sbox_1_and_788 ^ state_4_4_18_lpi_3
      ^ state_2_18_1_lpi_4 ^ state_1_1_31_0_lpi_4_18 ^ Encrypt_Top_sbox_1_and_798
      ^ state_4_4_23_lpi_3 ^ state_2_23_1_lpi_4 ^ state_1_1_31_0_lpi_4_23);
  assign xor_39_nl = state_2_17_1_lpi_4 ^ (key4[17]);
  assign state_xnor_16_nl = ~(xor_cse_483 ^ xor_cse_495 ^ state_4_3_31_0_sva_19 ^
      state_2_19_1_lpi_4 ^ plaintext_31_0_sva_19 ^ xor_cse_532 ^ state_4_3_31_0_sva_24
      ^ state_2_24_1_lpi_4 ^ plaintext_31_0_sva_24);
  assign state_xnor_17_nl = ~(Encrypt_Top_sbox_1_and_788 ^ state_4_4_18_lpi_3 ^ state_2_18_1_lpi_4
      ^ state_1_1_31_0_lpi_4_18 ^ Encrypt_Top_sbox_1_and_790 ^ state_4_4_19_lpi_3
      ^ state_2_19_1_lpi_4 ^ state_1_1_31_0_lpi_4_19 ^ Encrypt_Top_sbox_1_and_800
      ^ state_4_4_24_lpi_3 ^ state_2_24_1_lpi_4 ^ state_1_1_31_0_lpi_4_24);
  assign xor_37_nl = state_2_18_1_lpi_4 ^ (key4[18]);
  assign state_xnor_18_nl = ~(xor_cse_495 ^ state_4_3_31_0_sva_19 ^ state_2_19_1_lpi_4
      ^ plaintext_31_0_sva_19 ^ xor_cse_503 ^ state_4_3_31_0_sva_20 ^ state_2_20_1_lpi_4
      ^ plaintext_31_0_sva_20 ^ xor_cse_535 ^ state_4_3_31_0_sva_25 ^ state_2_25_1_lpi_4
      ^ plaintext_31_0_sva_25);
  assign state_xnor_19_nl = ~(Encrypt_Top_sbox_1_and_790 ^ state_4_4_19_lpi_3 ^ state_2_19_1_lpi_4
      ^ state_1_1_31_0_lpi_4_19 ^ Encrypt_Top_sbox_1_and_792 ^ state_4_4_20_lpi_3
      ^ state_2_20_1_lpi_4 ^ state_1_1_31_0_lpi_4_20 ^ Encrypt_Top_sbox_1_and_802
      ^ state_4_4_25_lpi_3 ^ state_2_25_1_lpi_4 ^ state_1_1_31_0_lpi_4_25);
  assign xor_35_nl = state_2_19_1_lpi_4 ^ (key4[19]);
  assign state_xnor_20_nl = ~(xor_cse_503 ^ state_4_3_31_0_sva_20 ^ state_2_20_1_lpi_4
      ^ plaintext_31_0_sva_20 ^ xor_cse_511 ^ state_4_3_31_0_sva_21 ^ state_2_21_1_lpi_4
      ^ plaintext_31_0_sva_21 ^ xor_cse_538 ^ state_4_3_31_0_sva_26 ^ state_2_26_1_lpi_4
      ^ plaintext_31_0_sva_26);
  assign state_xnor_21_nl = ~(xor_cse_539 ^ xor_cse_505 ^ xor_cse_513);
  assign xor_33_nl = state_2_20_1_lpi_4 ^ (key4[20]);
  assign state_xnor_22_nl = ~(xor_cse_511 ^ state_4_3_31_0_sva_21 ^ state_2_21_1_lpi_4
      ^ plaintext_31_0_sva_21 ^ xor_cse_519 ^ state_4_3_31_0_sva_22 ^ state_2_22_1_lpi_4
      ^ plaintext_31_0_sva_22 ^ xor_cse_543 ^ state_4_3_31_0_sva_27 ^ state_2_27_1_lpi_4
      ^ plaintext_31_0_sva_27);
  assign state_xnor_23_nl = ~(xor_cse_544 ^ xor_cse_513 ^ xor_cse_546);
  assign xor_31_nl = state_2_21_1_lpi_4 ^ (key4[21]);
  assign state_xnor_24_nl = ~(xor_cse_519 ^ state_4_3_31_0_sva_22 ^ state_2_22_1_lpi_4
      ^ plaintext_31_0_sva_22 ^ xor_cse_525 ^ state_4_3_31_0_sva_23 ^ state_2_23_1_lpi_4
      ^ plaintext_31_0_sva_23 ^ xor_cse_548 ^ state_4_3_31_0_sva_28 ^ state_2_28_1_lpi_4
      ^ plaintext_31_0_sva_28);
  assign state_xnor_25_nl = ~(xor_cse_549 ^ xor_cse_546 ^ xor_cse_551);
  assign xor_29_nl = state_2_22_1_lpi_4 ^ (key4[22]);
  assign state_xnor_26_nl = ~(xor_cse_525 ^ state_4_3_31_0_sva_23 ^ state_2_23_1_lpi_4
      ^ plaintext_31_0_sva_23 ^ xor_cse_532 ^ state_4_3_31_0_sva_24 ^ state_2_24_1_lpi_4
      ^ plaintext_31_0_sva_24 ^ xor_cse_553 ^ state_4_3_31_0_sva_29 ^ state_2_29_1_lpi_4
      ^ plaintext_31_0_sva_29);
  assign state_xnor_27_nl = ~(xor_cse_554 ^ xor_cse_551 ^ xor_cse_556);
  assign xor_27_nl = state_2_23_1_lpi_4 ^ (key4[23]);
  assign state_xnor_28_nl = ~(xor_cse_532 ^ state_4_3_31_0_sva_24 ^ state_2_24_1_lpi_4
      ^ plaintext_31_0_sva_24 ^ xor_cse_535 ^ state_4_3_31_0_sva_25 ^ state_2_25_1_lpi_4
      ^ plaintext_31_0_sva_25 ^ xor_cse_558 ^ state_4_3_31_0_sva_30 ^ state_2_30_1_lpi_4
      ^ plaintext_31_0_sva_30);
  assign state_xnor_29_nl = ~(xor_cse_559 ^ xor_cse_556 ^ xor_cse_561);
  assign xor_25_nl = state_2_24_1_lpi_4 ^ (key4[24]);
  assign state_xnor_30_nl = ~(xor_cse_535 ^ state_4_3_31_0_sva_25 ^ state_2_25_1_lpi_4
      ^ plaintext_31_0_sva_25 ^ xor_cse_538 ^ state_4_3_31_0_sva_26 ^ state_2_26_1_lpi_4
      ^ plaintext_31_0_sva_26 ^ xor_cse_565 ^ state_4_3_31_0_sva_31 ^ state_2_31_1_lpi_4
      ^ plaintext_31_0_sva_31);
  assign state_xnor_31_nl = ~(xor_cse_566 ^ xor_cse_539 ^ xor_cse_561);
  assign xor_23_nl = state_2_25_1_lpi_4 ^ (key4[25]);
  assign state_xnor_32_nl = ~(xor_cse_571 ^ xor_cse_538 ^ state_4_3_31_0_sva_26 ^
      state_2_26_1_lpi_4 ^ plaintext_31_0_sva_26 ^ xor_cse_574);
  assign state_xnor_33_nl = ~(xor_cse_544 ^ xor_cse_575 ^ xor_cse_539);
  assign xor_21_nl = state_2_26_1_lpi_4 ^ (key4[26]);
  assign state_xnor_34_nl = ~(xor_cse_544 ^ xor_cse_539 ^ xor_cse_576);
  assign state_xnor_35_nl = ~(xor_cse_581 ^ xor_cse_574 ^ xor_cse_548 ^ state_4_3_31_0_sva_28
      ^ state_2_28_1_lpi_4 ^ plaintext_31_0_sva_28);
  assign state_xnor_36_nl = ~(xor_cse_544 ^ xor_cse_585 ^ xor_cse_549);
  assign xor_19_nl = state_2_27_1_lpi_4 ^ (key4[27]);
  assign state_xnor_37_nl = ~(xor_cse_544 ^ xor_cse_549 ^ xor_cse_586);
  assign state_xnor_38_nl = ~(xor_cse_548 ^ state_4_3_31_0_sva_28 ^ state_2_28_1_lpi_4
      ^ plaintext_31_0_sva_28 ^ xor_cse_553 ^ state_4_3_31_0_sva_29 ^ state_2_29_1_lpi_4
      ^ plaintext_31_0_sva_29 ^ xor_cse_590 ^ state_4_3_63_32_sva_2 ^ state_2_34_1_lpi_4
      ^ plaintext_63_32_sva_2);
  assign state_xnor_39_nl = ~(xor_cse_591 ^ xor_cse_554 ^ state_4_4_28_lpi_3 ^ state_2_28_1_lpi_4
      ^ state_1_1_31_0_lpi_4_28 ^ state_1_1_63_32_lpi_4_2);
  assign xor_17_nl = state_2_28_1_lpi_4 ^ (key4[28]);
  assign state_xnor_40_nl = ~(xor_cse_591 ^ xor_cse_554 ^ state_4_4_28_lpi_3 ^ state_2_28_1_lpi_4
      ^ state_1_1_31_0_lpi_4_28 ^ state_1_1_63_32_lpi_4_0);
  assign state_xnor_41_nl = ~(xor_cse_597 ^ xor_cse_553 ^ state_4_3_31_0_sva_29 ^
      state_2_29_1_lpi_4 ^ plaintext_31_0_sva_29 ^ xor_cse_558 ^ state_4_3_31_0_sva_30
      ^ state_2_30_1_lpi_4 ^ plaintext_31_0_sva_30);
  assign state_xnor_42_nl = ~(xor_cse_559 ^ xor_cse_601 ^ xor_cse_554);
  assign xor_15_nl = state_2_29_1_lpi_4 ^ (key4[29]);
  assign state_xnor_43_nl = ~(xor_cse_559 ^ xor_cse_554 ^ xor_cse_602);
  assign state_xnor_44_nl = ~(xor_cse_558 ^ state_4_3_31_0_sva_30 ^ state_2_30_1_lpi_4
      ^ plaintext_31_0_sva_30 ^ xor_cse_565 ^ state_4_3_31_0_sva_31 ^ state_2_31_1_lpi_4
      ^ plaintext_31_0_sva_31 ^ xor_cse_606 ^ state_4_3_63_32_sva_4 ^ state_2_36_1_lpi_4
      ^ plaintext_63_32_sva_4);
  assign state_xnor_45_nl = ~(xor_cse_559 ^ xor_cse_566 ^ xor_cse_607);
  assign xor_13_nl = state_2_30_1_lpi_4 ^ (key4[30]);
  assign state_xnor_46_nl = ~(xor_cse_559 ^ xor_cse_608 ^ xor_cse_566);
  assign state_xnor_47_nl = ~(xor_cse_571 ^ xor_cse_565 ^ state_4_3_31_0_sva_31 ^
      state_2_31_1_lpi_4 ^ plaintext_31_0_sva_31 ^ xor_cse_613);
  assign state_xnor_48_nl = ~(xor_cse_575 ^ xor_cse_566 ^ Encrypt_Top_sbox_1_and_826
      ^ state_4_4_37_lpi_3 ^ state_2_37_1_lpi_4 ^ state_1_1_63_32_lpi_4_5);
  assign xor_7_nl = state_2_31_1_lpi_4 ^ (key4[31]);
  assign state_xnor_49_nl = ~(xor_cse_616 ^ xor_cse_566 ^ xor_cse_576);
  assign state_xnor_50_nl = ~(xor_cse_581 ^ xor_cse_571 ^ xor_cse_621);
  assign state_xnor_51_nl = ~(xor_cse_575 ^ xor_cse_585 ^ Encrypt_Top_sbox_1_and_828
      ^ state_4_4_38_lpi_3 ^ state_2_38_1_lpi_4 ^ state_1_1_63_32_lpi_4_6);
  assign state_xnor_52_nl = ~(xor_cse_624 ^ xor_cse_586 ^ xor_cse_576);
  assign state_xnor_53_nl = ~(xor_cse_581 ^ xor_cse_628 ^ xor_cse_629);
  assign state_xnor_54_nl = ~(xor_cse_585 ^ xor_cse_631 ^ Encrypt_Top_sbox_1_and_830
      ^ state_4_4_39_lpi_3 ^ state_2_39_1_lpi_4 ^ state_1_1_63_32_lpi_4_7);
  assign state_xnor_55_nl = ~(xor_cse_633 ^ xor_cse_586 ^ xor_cse_634);
  assign state_xnor_56_nl = ~(xor_cse_597 ^ xor_cse_637 ^ xor_cse_628);
  assign state_xnor_57_nl = ~(xor_cse_601 ^ xor_cse_631 ^ Encrypt_Top_sbox_1_and_832
      ^ state_4_4_40_lpi_3 ^ state_2_40_1_lpi_4 ^ state_1_1_63_32_lpi_4_8);
  assign state_xnor_58_nl = ~(xor_cse_641 ^ xor_cse_602 ^ xor_cse_634);
  assign state_xnor_59_nl = ~(xor_cse_597 ^ xor_cse_645 ^ xor_cse_606 ^ state_4_3_63_32_sva_4
      ^ state_2_36_1_lpi_4 ^ plaintext_63_32_sva_4);
  assign state_xnor_60_nl = ~(xor_cse_601 ^ xor_cse_607 ^ Encrypt_Top_sbox_1_and_834
      ^ state_4_4_41_lpi_3 ^ state_2_41_1_lpi_4 ^ state_1_1_63_32_lpi_4_9);
  assign state_xnor_61_nl = ~(xor_cse_650 ^ xor_cse_608 ^ xor_cse_602);
  assign state_xnor_62_nl = ~(xor_cse_606 ^ state_4_3_63_32_sva_4 ^ state_2_36_1_lpi_4
      ^ plaintext_63_32_sva_4 ^ xor_cse_614 ^ state_4_3_63_32_sva_5 ^ state_2_37_1_lpi_4
      ^ plaintext_63_32_sva_5 ^ xor_cse_653 ^ state_4_3_63_32_sva_10 ^ state_2_42_1_lpi_4
      ^ plaintext_63_32_sva_10);
  assign state_xnor_63_nl = ~(xor_cse_608 ^ state_1_1_63_32_lpi_4_4 ^ Encrypt_Top_sbox_1_and_826
      ^ state_4_4_37_lpi_3 ^ state_2_37_1_lpi_4 ^ state_1_1_63_32_lpi_4_5 ^ Encrypt_Top_sbox_1_and_836
      ^ state_4_4_42_lpi_3 ^ state_2_42_1_lpi_4);
  assign state_xnor_64_nl = ~(xor_cse_656 ^ xor_cse_616 ^ xor_cse_608);
  assign state_xnor_65_nl = ~(xor_cse_621 ^ xor_cse_659 ^ xor_cse_613);
  assign state_xnor_66_nl = ~(xor_cse_616 ^ state_1_1_63_32_lpi_4_5 ^ Encrypt_Top_sbox_1_and_828
      ^ state_4_4_38_lpi_3 ^ state_2_38_1_lpi_4 ^ state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_1_and_838
      ^ state_4_4_43_lpi_3 ^ state_2_43_1_lpi_4);
  assign state_xnor_67_nl = ~(xor_cse_624 ^ xor_cse_616 ^ xor_cse_664);
  assign state_xnor_68_nl = ~(xor_cse_621 ^ xor_cse_667 ^ xor_cse_629);
  assign state_xnor_69_nl = ~(xor_cse_624 ^ state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_1_and_830
      ^ state_4_4_39_lpi_3 ^ state_2_39_1_lpi_4 ^ state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_1_and_840
      ^ state_4_4_44_lpi_3 ^ state_2_44_1_lpi_4);
  assign state_xnor_70_nl = ~(xor_cse_624 ^ xor_cse_672 ^ xor_cse_633);
  assign state_xnor_71_nl = ~(xor_cse_637 ^ xor_cse_629 ^ xor_cse_676);
  assign state_xnor_72_nl = ~(xor_cse_633 ^ state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_1_and_832
      ^ state_4_4_40_lpi_3 ^ state_2_40_1_lpi_4 ^ state_1_1_63_32_lpi_4_8 ^ Encrypt_Top_sbox_1_and_842
      ^ state_4_4_45_lpi_3 ^ state_2_45_1_lpi_4);
  assign state_xnor_73_nl = ~(xor_cse_641 ^ xor_cse_633 ^ xor_cse_680);
  assign state_xnor_74_nl = ~(xor_cse_637 ^ xor_cse_645 ^ xor_cse_683);
  assign state_xnor_75_nl = ~(xor_cse_685 ^ state_1_1_63_32_lpi_4_9 ^ state_1_1_63_32_lpi_4_8
      ^ Encrypt_Top_sbox_1_and_834 ^ state_4_4_41_lpi_3 ^ state_2_41_1_lpi_4);
  assign state_xnor_76_nl = ~(state_1_1_63_32_lpi_4_2 ^ xor_cse_650 ^ xor_cse_685);
  assign state_xnor_77_nl = ~(xor_cse_645 ^ xor_cse_689 ^ xor_cse_690);
  assign state_xnor_78_nl = ~(xor_cse_650 ^ state_1_1_63_32_lpi_4_9 ^ Encrypt_Top_sbox_1_and_836
      ^ state_4_4_42_lpi_3 ^ state_2_42_1_lpi_4 ^ state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_1_and_846
      ^ state_4_4_47_lpi_3 ^ state_2_47_1_lpi_4);
  assign state_xnor_79_nl = ~(xor_cse_656 ^ xor_cse_650 ^ xor_cse_694);
  assign state_xnor_80_nl = ~(xor_cse_659 ^ xor_cse_689 ^ xor_cse_698 ^ state_4_3_63_32_sva_16
      ^ state_2_48_1_lpi_4 ^ plaintext_63_32_sva_16);
  assign state_xnor_81_nl = ~(xor_cse_656 ^ state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_1_and_838
      ^ state_4_4_43_lpi_3 ^ state_2_43_1_lpi_4 ^ state_1_1_63_32_lpi_4_11 ^ Encrypt_Top_sbox_1_and_848
      ^ state_4_4_48_lpi_3 ^ state_2_48_1_lpi_4);
  assign state_xnor_82_nl = ~(xor_cse_656 ^ xor_cse_701 ^ xor_cse_664);
  assign state_xnor_83_nl = ~(xor_cse_659 ^ xor_cse_667 ^ xor_cse_705 ^ state_4_3_63_32_sva_17
      ^ state_2_49_1_lpi_4 ^ plaintext_63_32_sva_17);
  assign state_xnor_84_nl = ~(xor_cse_664 ^ state_1_1_63_32_lpi_4_11 ^ Encrypt_Top_sbox_1_and_840
      ^ state_4_4_44_lpi_3 ^ state_2_44_1_lpi_4 ^ state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_1_and_850
      ^ state_4_4_49_lpi_3 ^ state_2_49_1_lpi_4);
  assign state_xnor_85_nl = ~(xor_cse_708 ^ xor_cse_672 ^ xor_cse_664);
  assign state_xnor_86_nl = ~(xor_cse_667 ^ xor_cse_676 ^ xor_cse_713 ^ state_4_3_63_32_sva_18
      ^ state_2_50_1_lpi_4 ^ plaintext_63_32_sva_18);
  assign state_xnor_87_nl = ~(xor_cse_672 ^ state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_1_and_842
      ^ state_4_4_45_lpi_3 ^ state_2_45_1_lpi_4 ^ state_1_1_63_32_lpi_4_13 ^ Encrypt_Top_sbox_1_and_852
      ^ state_4_4_50_lpi_3 ^ state_2_50_1_lpi_4);
  assign state_xnor_88_nl = ~(xor_cse_672 ^ xor_cse_716 ^ xor_cse_680);
  assign state_xnor_89_nl = ~(xor_cse_683 ^ xor_cse_676 ^ xor_cse_721 ^ state_4_3_63_32_sva_19
      ^ state_2_51_1_lpi_4 ^ plaintext_63_32_sva_19);
  assign state_xnor_90_nl = ~(xor_cse_680 ^ xor_cse_722 ^ state_1_1_63_32_lpi_4_13
      ^ Encrypt_Top_sbox_1_and_854 ^ state_4_4_51_lpi_3 ^ state_2_51_1_lpi_4);
  assign state_xnor_91_nl = ~(xor_cse_724 ^ xor_cse_680 ^ xor_cse_725);
  assign state_xnor_92_nl = ~(xor_cse_683 ^ xor_cse_690 ^ xor_cse_730 ^ state_4_3_63_32_sva_20
      ^ state_2_52_1_lpi_4 ^ plaintext_63_32_sva_20);
  assign state_xnor_93_nl = ~(xor_cse_694 ^ xor_cse_722 ^ state_1_1_63_32_lpi_4_15
      ^ Encrypt_Top_sbox_1_and_856 ^ state_4_4_52_lpi_3 ^ state_2_52_1_lpi_4);
  assign state_xnor_94_nl = ~(xor_cse_732 ^ xor_cse_694 ^ xor_cse_725);
  assign state_xnor_95_nl = ~(xor_cse_691 ^ state_4_3_63_32_sva_15 ^ state_2_47_1_lpi_4
      ^ plaintext_63_32_sva_15 ^ xor_cse_698 ^ state_4_3_63_32_sva_16 ^ state_2_48_1_lpi_4
      ^ plaintext_63_32_sva_16 ^ xor_cse_736 ^ state_4_3_63_32_sva_21 ^ state_2_53_1_lpi_4
      ^ plaintext_63_32_sva_21);
  assign state_xnor_96_nl = ~(xor_cse_701 ^ Encrypt_Top_sbox_1_and_846 ^ state_4_4_47_lpi_3
      ^ state_2_47_1_lpi_4 ^ state_1_1_63_32_lpi_4_15 ^ state_1_1_63_32_lpi_4_16
      ^ Encrypt_Top_sbox_1_and_858 ^ state_4_4_53_lpi_3 ^ state_2_53_1_lpi_4);
  assign state_xnor_97_nl = ~(xor_cse_739 ^ xor_cse_694 ^ xor_cse_701);
  assign state_xnor_98_nl = ~(xor_cse_698 ^ state_4_3_63_32_sva_16 ^ state_2_48_1_lpi_4
      ^ plaintext_63_32_sva_16 ^ xor_cse_705 ^ state_4_3_63_32_sva_17 ^ state_2_49_1_lpi_4
      ^ plaintext_63_32_sva_17 ^ xor_cse_742 ^ state_4_3_63_32_sva_22 ^ state_2_54_1_lpi_4
      ^ plaintext_63_32_sva_22);
  assign state_xnor_99_nl = ~(xor_cse_743 ^ state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_1_and_848
      ^ state_4_4_48_lpi_3 ^ state_2_48_1_lpi_4 ^ state_1_1_63_32_lpi_4_16);
  assign state_xnor_100_nl = ~(state_1_1_63_32_lpi_4_27 ^ xor_cse_701 ^ xor_cse_743);
  assign state_xnor_101_nl = ~(xor_cse_705 ^ state_4_3_63_32_sva_17 ^ state_2_49_1_lpi_4
      ^ plaintext_63_32_sva_17 ^ xor_cse_713 ^ state_4_3_63_32_sva_18 ^ state_2_50_1_lpi_4
      ^ plaintext_63_32_sva_18 ^ xor_cse_748 ^ state_4_3_63_32_sva_23 ^ state_2_55_1_lpi_4
      ^ plaintext_63_32_sva_23);
  assign state_xnor_102_nl = ~(xor_cse_749 ^ state_1_1_63_32_lpi_4_18 ^ Encrypt_Top_sbox_1_and_850
      ^ state_4_4_49_lpi_3 ^ state_2_49_1_lpi_4 ^ state_1_1_63_32_lpi_4_17);
  assign state_xnor_103_nl = ~(state_1_1_63_32_lpi_4_28 ^ xor_cse_708 ^ xor_cse_749);
  assign state_xnor_104_nl = ~(xor_cse_713 ^ state_4_3_63_32_sva_18 ^ state_2_50_1_lpi_4
      ^ plaintext_63_32_sva_18 ^ xor_cse_721 ^ state_4_3_63_32_sva_19 ^ state_2_51_1_lpi_4
      ^ plaintext_63_32_sva_19 ^ xor_cse_754 ^ state_4_3_63_32_sva_24 ^ state_2_56_1_lpi_4
      ^ plaintext_63_32_sva_24);
  assign state_xnor_105_nl = ~(xor_cse_755 ^ state_1_1_63_32_lpi_4_19 ^ Encrypt_Top_sbox_1_and_852
      ^ state_4_4_50_lpi_3 ^ state_2_50_1_lpi_4 ^ state_1_1_63_32_lpi_4_18);
  assign state_xnor_106_nl = ~(state_1_1_63_32_lpi_4_29 ^ xor_cse_716 ^ xor_cse_755);
  assign state_xnor_107_nl = ~(xor_cse_721 ^ state_4_3_63_32_sva_19 ^ state_2_51_1_lpi_4
      ^ plaintext_63_32_sva_19 ^ xor_cse_730 ^ state_4_3_63_32_sva_20 ^ state_2_52_1_lpi_4
      ^ plaintext_63_32_sva_20 ^ xor_cse_759 ^ state_4_3_63_32_sva_25 ^ state_2_57_1_lpi_4
      ^ plaintext_63_32_sva_25);
  assign state_xnor_108_nl = ~(xor_cse_760 ^ state_1_1_63_32_lpi_4_20 ^ Encrypt_Top_sbox_1_and_854
      ^ state_4_4_51_lpi_3 ^ state_2_51_1_lpi_4 ^ state_1_1_63_32_lpi_4_19);
  assign state_xnor_109_nl = ~(state_1_1_63_32_lpi_4_3 ^ xor_cse_724 ^ xor_cse_760);
  assign state_xnor_110_nl = ~(xor_cse_730 ^ state_4_3_63_32_sva_20 ^ state_2_52_1_lpi_4
      ^ plaintext_63_32_sva_20 ^ xor_cse_736 ^ state_4_3_63_32_sva_21 ^ state_2_53_1_lpi_4
      ^ plaintext_63_32_sva_21 ^ xor_cse_764 ^ state_4_3_63_32_sva_26 ^ state_2_58_1_lpi_4
      ^ plaintext_63_32_sva_26);
  assign state_xnor_111_nl = ~(xor_cse_739 ^ Encrypt_Top_sbox_1_and_868 ^ Encrypt_Top_sbox_1_and_856
      ^ state_4_4_52_lpi_3 ^ state_2_52_1_lpi_4 ^ state_1_1_63_32_lpi_4_20 ^ state_1_1_63_32_lpi_4_21
      ^ state_4_4_58_lpi_3 ^ state_2_58_1_lpi_4);
  assign state_xnor_112_nl = ~(xor_cse_739 ^ xor_cse_732 ^ xor_cse_767);
  assign state_xnor_113_nl = ~(xor_cse_736 ^ state_4_3_63_32_sva_21 ^ state_2_53_1_lpi_4
      ^ plaintext_63_32_sva_21 ^ xor_cse_742 ^ state_4_3_63_32_sva_22 ^ state_2_54_1_lpi_4
      ^ plaintext_63_32_sva_22 ^ xor_cse_769 ^ state_4_3_63_32_sva_27 ^ state_2_59_1_lpi_4
      ^ plaintext_63_32_sva_27);
  assign state_xnor_114_nl = ~(xor_cse_770 ^ xor_cse_771 ^ Encrypt_Top_sbox_1_and_858
      ^ state_4_4_53_lpi_3 ^ state_2_53_1_lpi_4 ^ state_1_1_63_32_lpi_4_21);
  assign state_xnor_115_nl = ~(xor_cse_770 ^ xor_cse_739 ^ Encrypt_Top_sbox_1_and_860
      ^ state_4_4_54_lpi_3 ^ state_2_54_1_lpi_4 ^ state_1_1_63_32_lpi_4_31);
  assign state_xnor_116_nl = ~(xor_cse_742 ^ state_4_3_63_32_sva_22 ^ state_2_54_1_lpi_4
      ^ plaintext_63_32_sva_22 ^ xor_cse_748 ^ state_4_3_63_32_sva_23 ^ state_2_55_1_lpi_4
      ^ plaintext_63_32_sva_23 ^ xor_cse_776 ^ state_4_3_63_32_sva_28 ^ state_2_60_1_lpi_4
      ^ plaintext_63_32_sva_28);
  assign state_xnor_117_nl = ~(xor_cse_777 ^ xor_cse_771 ^ Encrypt_Top_sbox_1_and_862
      ^ state_4_4_55_lpi_3 ^ state_2_55_1_lpi_4 ^ state_1_1_63_32_lpi_4_23);
  assign state_xnor_118_nl = ~(xor_cse_777 ^ Encrypt_Top_sbox_1_and_860 ^ state_4_4_54_lpi_3
      ^ state_2_54_1_lpi_4 ^ state_1_1_63_32_lpi_4_27 ^ Encrypt_Top_sbox_1_and_862
      ^ state_4_4_55_lpi_3 ^ state_2_55_1_lpi_4 ^ state_1_1_63_32_lpi_4_4);
  assign state_xnor_119_nl = ~(xor_cse_748 ^ state_4_3_63_32_sva_23 ^ state_2_55_1_lpi_4
      ^ plaintext_63_32_sva_23 ^ xor_cse_754 ^ state_4_3_63_32_sva_24 ^ state_2_56_1_lpi_4
      ^ plaintext_63_32_sva_24 ^ xor_cse_782 ^ state_4_3_63_32_sva_29 ^ state_2_61_1_lpi_4
      ^ plaintext_63_32_sva_29);
  assign state_xnor_120_nl = ~(xor_cse_783 ^ xor_cse_784 ^ state_1_1_63_32_lpi_4_23
      ^ state_4_4_56_lpi_3 ^ state_2_56_1_lpi_4 ^ state_1_1_63_32_lpi_4_24);
  assign state_xnor_121_nl = ~(xor_cse_783 ^ xor_cse_784 ^ state_1_1_63_32_lpi_4_28
      ^ state_4_4_56_lpi_3 ^ state_2_56_1_lpi_4 ^ state_1_1_63_32_lpi_4_5);
  assign state_xnor_122_nl = ~(xor_cse_754 ^ state_4_3_63_32_sva_24 ^ state_2_56_1_lpi_4
      ^ plaintext_63_32_sva_24 ^ xor_cse_759 ^ state_4_3_63_32_sva_25 ^ state_2_57_1_lpi_4
      ^ plaintext_63_32_sva_25 ^ xor_cse_788 ^ state_4_3_63_32_sva_30 ^ state_2_62_1_lpi_4
      ^ plaintext_63_32_sva_30);
  assign state_xnor_123_nl = ~(xor_cse_789 ^ xor_cse_790 ^ state_1_1_63_32_lpi_4_24
      ^ state_4_4_57_lpi_3 ^ state_2_57_1_lpi_4 ^ state_1_1_63_32_lpi_4_25);
  assign state_xnor_124_nl = ~(xor_cse_790 ^ xor_cse_792 ^ state_1_1_63_32_lpi_4_29
      ^ state_4_4_57_lpi_3 ^ state_2_57_1_lpi_4 ^ state_1_1_63_32_lpi_4_3);
  assign state_xnor_125_nl = ~(xor_cse_759 ^ state_4_3_63_32_sva_25 ^ state_2_57_1_lpi_4
      ^ plaintext_63_32_sva_25 ^ xor_cse_764 ^ state_4_3_63_32_sva_26 ^ state_2_58_1_lpi_4
      ^ plaintext_63_32_sva_26 ^ xor_cse_795 ^ state_4_3_63_32_sva_31 ^ state_2_63_1_lpi_4
      ^ plaintext_63_32_sva_31);
  assign state_xnor_126_nl = ~(xor_cse_796 ^ xor_cse_797 ^ Encrypt_Top_sbox_1_and_866
      ^ state_4_4_57_lpi_3 ^ state_2_57_1_lpi_4 ^ state_1_1_63_32_lpi_4_25);
  assign state_xnor_127_nl = ~(xor_cse_767 ^ xor_cse_799 ^ Encrypt_Top_sbox_1_and_866
      ^ state_4_4_57_lpi_3 ^ state_2_57_1_lpi_4 ^ state_1_1_63_32_lpi_4_3);
  assign state_xnor_146_nl = ~(xor_cse_845 ^ xor_cse_847 ^ xor_cse_494 ^ state_4_3_31_0_sva_14
      ^ state_2_14_1_lpi_4 ^ plaintext_31_0_sva_14);
  assign state_xnor_147_nl = ~(xor_cse_850 ^ xor_cse_851 ^ xor_cse_496);
  assign state_xnor_148_nl = ~(xor_cse_852 ^ xor_cse_496 ^ Encrypt_Top_sbox_1_and_880
      ^ state_4_4_8_lpi_3 ^ state_2_8_1_lpi_4 ^ state_1_1_63_32_lpi_4_8);
  assign state_xnor_149_nl = ~(xor_cse_847 ^ xor_cse_461 ^ xor_cse_509);
  assign state_xnor_150_nl = ~(xor_cse_465 ^ xor_cse_504 ^ xor_cse_851);
  assign state_xnor_151_nl = ~(xor_cse_465 ^ xor_cse_852 ^ xor_cse_504);
  assign state_xnor_128_nl = ~(plaintext_31_0_sva_0 ^ xor_cse_802 ^ xor_cse_764 ^
      state_4_3_63_32_sva_26 ^ state_2_58_1_lpi_4 ^ plaintext_63_32_sva_26 ^ xor_cse_805);
  assign state_xnor_129_nl = ~(state_2_0_1_lpi_4 ^ xor_cse_770 ^ xor_cse_806 ^ xor_cse_797);
  assign Encrypt_Top_linear_2_xnor_nl = ~(state_2_0_1_lpi_6 ^ xor_cse_770 ^ xor_cse_806
      ^ xor_cse_797);
  assign xor_64_nl = state_2_58_1_lpi_4 ^ (key3[26]);
  assign state_xnor_130_nl = ~(state_1_1_31_0_lpi_4_0 ^ xor_cse_767 ^ xor_cse_807
      ^ xor_cse_808);
  assign state_xnor_131_nl = ~(plaintext_31_0_sva_1 ^ xor_cse_809 ^ xor_cse_805 ^
      xor_cse_812);
  assign state_xnor_132_nl = ~(state_2_1_1_lpi_4 ^ xor_cse_777 ^ xor_cse_770 ^ xor_cse_813);
  assign Encrypt_Top_linear_2_xnor_1_nl = ~(state_2_1_1_lpi_6 ^ xor_cse_777 ^ xor_cse_770
      ^ xor_cse_813);
  assign xor_66_nl = state_2_59_1_lpi_4 ^ (key3[27]);
  assign state_xnor_133_nl = ~(state_1_1_31_0_lpi_4_1 ^ xor_cse_814 ^ xor_cse_807
      ^ Encrypt_Top_sbox_1_and_872 ^ state_4_4_60_lpi_3 ^ state_2_60_1_lpi_4 ^ state_1_1_63_32_lpi_4_4);
  assign state_xnor_134_nl = ~(plaintext_31_0_sva_2 ^ xor_cse_817 ^ xor_cse_812 ^
      xor_cse_820);
  assign state_xnor_135_nl = ~(state_2_2_1_lpi_4 ^ xor_cse_783 ^ xor_cse_777 ^ xor_cse_821);
  assign Encrypt_Top_linear_2_xnor_2_nl = ~(state_2_2_1_lpi_6 ^ xor_cse_783 ^ xor_cse_777
      ^ xor_cse_821);
  assign xor_68_nl = state_2_60_1_lpi_4 ^ (key3[28]);
  assign state_xnor_136_nl = ~(Encrypt_Top_sbox_1_and_872 ^ state_4_4_60_lpi_3 ^
      state_2_60_1_lpi_4 ^ state_1_1_63_32_lpi_4_4 ^ Encrypt_Top_sbox_1_and_874 ^
      state_4_4_61_lpi_3 ^ state_2_61_1_lpi_4 ^ state_1_1_63_32_lpi_4_5 ^ Encrypt_Top_sbox_1_and_760
      ^ state_4_4_2_lpi_3 ^ state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ state_1_1_31_0_lpi_4_2);
  assign state_xnor_137_nl = ~(plaintext_31_0_sva_3 ^ xor_cse_822 ^ xor_cse_820 ^
      xor_cse_825);
  assign state_xnor_138_nl = ~(state_2_3_1_lpi_4 ^ xor_cse_783 ^ xor_cse_789 ^ xor_cse_826);
  assign Encrypt_Top_linear_2_xnor_3_nl = ~(state_2_3_1_lpi_6 ^ xor_cse_783 ^ xor_cse_789
      ^ xor_cse_826);
  assign xor_70_nl = state_2_61_1_lpi_4 ^ (key3[29]);
  assign state_xnor_139_nl = ~(state_1_1_31_0_lpi_4_3 ^ xor_cse_792 ^ xor_cse_827
      ^ Encrypt_Top_sbox_1_and_874 ^ state_4_4_61_lpi_3 ^ state_2_61_1_lpi_4 ^ state_1_1_63_32_lpi_4_5);
  assign state_xnor_140_nl = ~(plaintext_31_0_sva_4 ^ xor_cse_829 ^ xor_cse_825 ^
      xor_cse_832);
  assign state_xnor_141_nl = ~(state_2_4_1_lpi_4 ^ xor_cse_789 ^ xor_cse_796 ^ xor_cse_833);
  assign Encrypt_Top_linear_2_xnor_4_nl = ~(state_2_4_1_lpi_6 ^ xor_cse_789 ^ xor_cse_796
      ^ xor_cse_833);
  assign xor_72_nl = state_2_62_1_lpi_4 ^ (key3[30]);
  assign state_xnor_142_nl = ~(state_1_1_31_0_lpi_4_4 ^ xor_cse_834 ^ xor_cse_792
      ^ xor_cse_799);
  assign state_xnor_143_nl = ~(xor_cse_802 ^ xor_cse_835 ^ xor_cse_832 ^ plaintext_31_0_sva_0
      ^ plaintext_31_0_sva_5);
  assign state_xnor_144_nl = ~(xor_cse_796 ^ xor_cse_806 ^ xor_cse_839 ^ state_2_0_1_lpi_4
      ^ state_2_5_1_lpi_4);
  assign Encrypt_Top_linear_2_xnor_5_nl = ~(xor_cse_796 ^ xor_cse_806 ^ xor_cse_839
      ^ state_2_0_1_lpi_6 ^ state_2_5_1_lpi_6);
  assign xor_74_nl = state_2_63_1_lpi_4 ^ (key3[31]);
  assign state_xnor_145_nl = ~(xor_cse_842 ^ xor_cse_799 ^ xor_cse_808 ^ state_1_1_31_0_lpi_4_0
      ^ state_1_1_31_0_lpi_4_5);
  assign state_xor_82_nl = xor_cse_858 ^ xor_cse_366 ^ xor_cse_861 ^ Encrypt_Top_sbox_and_1_cse_10_sva_1
      ^ state_2_10_1_lpi_4 ^ state_0_10_lpi_6 ^ Encrypt_Top_sbox_and_1_cse_29_sva_1
      ^ state_2_29_1_lpi_4 ^ state_0_29_lpi_6;
  assign state_xor_83_nl = xor_cse_368 ^ xor_cse_272 ^ xor_cse_87 ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1
      ^ state_2_38_1_lpi_4 ^ state_0_38_lpi_6;
  assign state_xor_84_nl = xor_cse_368 ^ xor_cse_272 ^ xor_cse_866;
  assign mux1h_64_nl = MUX1HOT_s_1_5_2(state_xor_82_nl, state_0_10_sva_2_mx0w1, state_xor_83_nl,
      data_out_rsci_idat_10, state_xor_84_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_85_nl = Encrypt_Top_sbox_and_2_cse_39_sva_1 ^ xor_cse_867 ^ xor_cse_379
      ^ xor_cse_868 ^ Encrypt_Top_sbox_and_1_cse_11_sva_1 ^ state_2_11_1_lpi_4 ^
      state_0_11_lpi_6 ^ Encrypt_Top_sbox_and_1_cse_30_sva_1 ^ state_2_30_1_lpi_4
      ^ state_0_30_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_7 ^ Encrypt_Top_sbox_and_1_cse_39_sva_1;
  assign state_xor_86_nl = xor_cse_280 ^ xor_cse_871 ^ xor_cse_98 ^ Encrypt_Top_sbox_1_and_1_cse_39_sva_1
      ^ state_2_39_1_lpi_4 ^ state_0_39_lpi_6;
  assign state_xor_87_nl = xor_cse_280 ^ xor_cse_871 ^ xor_cse_875 ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1 ^ state_0_39_lpi_6;
  assign mux1h_65_nl = MUX1HOT_s_1_5_2(state_xor_85_nl, state_0_11_sva_2_mx0w1, state_xor_86_nl,
      data_out_rsci_idat_11, state_xor_87_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_88_nl = xor_cse_877 ^ xor_cse_390 ^ xor_cse_880 ^ Encrypt_Top_sbox_and_1_cse_12_sva_1
      ^ state_2_12_1_lpi_4 ^ state_0_12_lpi_6 ^ Encrypt_Top_sbox_and_1_cse_31_sva_1
      ^ state_2_31_1_lpi_4 ^ state_0_31_lpi_6;
  assign state_xor_89_nl = xor_cse_393 ^ xor_cse_288 ^ xor_cse_113 ^ Encrypt_Top_sbox_1_and_1_cse_40_sva_1
      ^ state_2_40_1_lpi_4 ^ state_0_40_lpi_6;
  assign state_xor_90_nl = xor_cse_393 ^ xor_cse_288 ^ xor_cse_635 ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1
      ^ state_2_40_1_lpi_4 ^ state_0_40_lpi_6;
  assign mux1h_66_nl = MUX1HOT_s_1_5_2(state_xor_88_nl, state_0_12_sva_2_mx0w1, state_xor_89_nl,
      data_out_rsci_idat_12, state_xor_90_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_91_nl = xor_cse_887 ^ xor_cse_400 ^ xor_cse_890 ^ Encrypt_Top_sbox_and_1_cse_13_sva_1
      ^ state_2_13_1_lpi_4 ^ state_0_13_lpi_6;
  assign state_xor_92_nl = xor_cse_297 ^ xor_cse_4 ^ xor_cse_128 ^ Encrypt_Top_sbox_1_and_1_cse_32_sva_1
      ^ state_2_32_1_lpi_4 ^ state_0_32_lpi_6 ^ Encrypt_Top_sbox_1_and_cse_41_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1 ^ state_0_41_lpi_6;
  assign state_xor_93_nl = xor_cse_297 ^ xor_cse_895 ^ xor_cse_897 ^ Encrypt_Top_sbox_3_and_1_cse_41_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_41_sva_1 ^ state_0_41_lpi_6;
  assign mux1h_67_nl = MUX1HOT_s_1_5_2(state_xor_91_nl, state_0_13_sva_2_mx0w1, state_xor_92_nl,
      data_out_rsci_idat_13, state_xor_93_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_94_nl = Encrypt_Top_sbox_and_2_cse_42_sva_1 ^ xor_cse_899 ^ xor_cse_419
      ^ xor_cse_900 ^ Encrypt_Top_sbox_and_1_cse_14_sva_1 ^ state_2_14_1_lpi_4 ^
      state_0_14_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_1 ^ Encrypt_Top_sbox_and_1_cse_33_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_33_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_10
      ^ Encrypt_Top_sbox_and_1_cse_42_sva_1;
  assign state_xor_95_nl = xor_cse_306 ^ xor_cse_140 ^ xor_cse_18 ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1
      ^ state_2_33_1_lpi_4 ^ state_0_33_lpi_6 ^ Encrypt_Top_sbox_1_and_cse_42_sva_1
      ^ xor_cse_905;
  assign state_xor_96_nl = xor_cse_306 ^ xor_cse_906 ^ xor_cse_651 ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1
      ^ state_2_42_1_lpi_4 ^ state_0_42_lpi_6;
  assign mux1h_68_nl = MUX1HOT_s_1_5_2(state_xor_94_nl, state_0_14_sva_2_mx0w1, state_xor_95_nl,
      data_out_rsci_idat_14, state_xor_96_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_97_nl = xor_cse_909 ^ xor_cse_431 ^ xor_cse_912 ^ Encrypt_Top_sbox_and_1_cse_15_sva_1
      ^ state_2_15_1_lpi_4 ^ state_0_15_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_2
      ^ Encrypt_Top_sbox_and_1_cse_34_sva_1 ^ Encrypt_Top_sbox_and_2_cse_34_sva_1;
  assign state_xor_98_nl = xor_cse_915 ^ xor_cse_231 ^ xor_cse_30 ^ state_0_34_lpi_6
      ^ Encrypt_Top_sbox_1_and_cse_15_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_15_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1
      ^ state_2_34_1_lpi_4;
  assign state_xor_99_nl = xor_cse_438 ^ xor_cse_231 ^ xor_cse_920 ^ Encrypt_Top_sbox_1_and_cse_15_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_15_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1
      ^ state_0_43_lpi_6;
  assign mux1h_69_nl = MUX1HOT_s_1_5_2(state_xor_97_nl, state_0_15_sva_2_mx0w1, state_xor_98_nl,
      data_out_rsci_idat_15, state_xor_99_nl, {(fsm_output[1]) , (fsm_output[3])
      , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_100_nl = xor_cse_445 ^ xor_cse_923 ^ xor_cse_926 ^ xor_cse_927;
  assign state_xor_101_nl = Encrypt_Top_sbox_2_and_2_cse_44_sva_1 ^ xor_cse_242 ^
      xor_cse_46 ^ xor_cse_160 ^ xor_cse_928 ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_35_sva_1 ^ state_2_35_1_lpi_4 ^ state_0_35_lpi_6;
  assign state_xor_102_nl = xor_cse_457 ^ xor_cse_242 ^ xor_cse_568 ^ xor_cse_928
      ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1;
  assign mux1h_70_nl = MUX1HOT_s_1_5_2(state_xor_100_nl, state_0_16_sva_2_mx0w1,
      state_xor_101_nl, data_out_rsci_idat_16, state_xor_102_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_103_nl = xor_cse_932 ^ xor_cse_935 ^ xor_cse_936 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_4
      ^ Encrypt_Top_sbox_and_1_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_36_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_13 ^ Encrypt_Top_sbox_and_1_cse_45_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_45_sva_1;
  assign state_xor_104_nl = xor_cse_251 ^ xor_cse_168 ^ xor_cse_59 ^ Encrypt_Top_sbox_1_and_1_cse_36_sva_1
      ^ state_2_36_1_lpi_4 ^ state_0_36_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_45_sva_1
      ^ state_2_45_1_lpi_4 ^ state_0_45_lpi_6;
  assign state_xor_105_nl = xor_cse_251 ^ xor_cse_943 ^ xor_cse_944 ^ Encrypt_Top_sbox_3_and_1_cse_36_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1 ^ state_0_36_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1 ^ state_0_45_lpi_6;
  assign mux1h_71_nl = MUX1HOT_s_1_5_2(state_xor_103_nl, state_0_17_sva_2_mx0w1,
      state_xor_104_nl, data_out_rsci_idat_17, state_xor_105_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_106_nl = xor_cse_947 ^ xor_cse_950 ^ xor_cse_951 ^ Encrypt_Top_sbox_and_1_cse_18_sva_1
      ^ state_2_18_1_lpi_4 ^ state_0_18_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_5
      ^ xor_cse_953;
  assign state_xor_107_nl = xor_cse_341 ^ xor_cse_181 ^ xor_cse_74 ^ xor_cse_955
      ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1 ^ state_2_37_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_46_sva_1;
  assign state_xor_108_nl = xor_cse_341 ^ xor_cse_958 ^ xor_cse_604 ^ xor_cse_955
      ^ Encrypt_Top_sbox_3_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_46_sva_1;
  assign mux1h_72_nl = MUX1HOT_s_1_5_2(state_xor_106_nl, state_0_18_sva_2_mx0w1,
      state_xor_107_nl, data_out_rsci_idat_18, state_xor_108_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_109_nl = xor_cse_349 ^ xor_cse_858 ^ xor_cse_961 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_15
      ^ Encrypt_Top_sbox_and_1_cse_47_sva_1 ^ Encrypt_Top_sbox_and_2_cse_47_sva_1;
  assign state_xor_110_nl = xor_cse_358 ^ xor_cse_192 ^ xor_cse_87 ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1
      ^ state_2_38_1_lpi_4 ^ state_0_38_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_47_sva_1
      ^ state_2_47_1_lpi_4 ^ state_0_47_lpi_6;
  assign state_xor_111_nl = xor_cse_358 ^ xor_cse_866 ^ xor_cse_967 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1 ^ state_0_47_lpi_6;
  assign mux1h_73_nl = MUX1HOT_s_1_5_2(state_xor_109_nl, state_0_19_sva_2_mx0w1,
      state_xor_110_nl, data_out_rsci_idat_19, state_xor_111_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_112_nl = xor_cse_361 ^ xor_cse_970 ^ xor_cse_867 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_7
      ^ Encrypt_Top_sbox_and_1_cse_39_sva_1 ^ Encrypt_Top_sbox_and_2_cse_39_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_16 ^ Encrypt_Top_sbox_and_1_cse_48_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_48_sva_1;
  assign state_xor_113_nl = xor_cse_370 ^ xor_cse_201 ^ xor_cse_98 ^ Encrypt_Top_sbox_1_and_1_cse_39_sva_1
      ^ state_2_39_1_lpi_4 ^ state_0_39_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_48_sva_1
      ^ state_2_48_1_lpi_4 ^ state_0_48_lpi_6;
  assign state_xor_114_nl = xor_cse_370 ^ xor_cse_875 ^ xor_cse_977 ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1 ^ state_0_39_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1 ^ state_0_48_lpi_6;
  assign mux1h_74_nl = MUX1HOT_s_1_5_2(state_xor_112_nl, state_0_20_sva_2_mx0w1,
      state_xor_113_nl, data_out_rsci_idat_20, state_xor_114_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_115_nl = xor_cse_374 ^ xor_cse_877 ^ xor_cse_981 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_17
      ^ Encrypt_Top_sbox_and_1_cse_49_sva_1 ^ Encrypt_Top_sbox_and_2_cse_49_sva_1;
  assign state_xor_116_nl = xor_cse_983 ^ xor_cse_214 ^ xor_cse_113 ^ xor_cse_985
      ^ Encrypt_Top_sbox_1_and_1_cse_40_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_49_sva_1;
  assign state_xor_117_nl = xor_cse_983 ^ xor_cse_702 ^ xor_cse_635 ^ xor_cse_985
      ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1;
  assign mux1h_75_nl = MUX1HOT_s_1_5_2(state_xor_115_nl, state_0_21_sva_2_mx0w1,
      state_xor_116_nl, data_out_rsci_idat_21, state_xor_117_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_118_nl = xor_cse_386 ^ xor_cse_887 ^ xor_cse_990 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_18
      ^ Encrypt_Top_sbox_and_1_cse_50_sva_1 ^ Encrypt_Top_sbox_and_2_cse_50_sva_1;
  assign state_xor_119_nl = xor_cse_395 ^ xor_cse_224 ^ xor_cse_128 ^ Encrypt_Top_sbox_1_and_cse_41_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1 ^ state_0_41_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_50_sva_1
      ^ state_2_50_1_lpi_4 ^ state_0_50_lpi_6;
  assign state_xor_120_nl = xor_cse_395 ^ xor_cse_897 ^ xor_cse_996 ^ Encrypt_Top_sbox_3_and_1_cse_41_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_41_sva_1 ^ state_0_41_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_50_sva_1 ^ state_0_50_lpi_6;
  assign mux1h_76_nl = MUX1HOT_s_1_5_2(state_xor_118_nl, state_0_22_sva_2_mx0w1,
      state_xor_119_nl, data_out_rsci_idat_22, state_xor_120_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_121_nl = xor_cse_402 ^ xor_cse_1000 ^ xor_cse_899 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_10
      ^ Encrypt_Top_sbox_and_1_cse_42_sva_1 ^ Encrypt_Top_sbox_and_2_cse_42_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_19 ^ Encrypt_Top_sbox_and_1_cse_51_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_51_sva_1;
  assign state_xor_122_nl = xor_cse ^ xor_cse_308 ^ xor_cse_140 ^ Encrypt_Top_sbox_1_and_cse_23_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_23_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1
      ^ Encrypt_Top_sbox_1_and_cse_42_sva_1 ^ xor_cse_905;
  assign state_xor_123_nl = state_0_51_lpi_6 ^ xor_cse_308 ^ xor_cse_651 ^ xor_cse_717
      ^ Encrypt_Top_sbox_1_and_cse_23_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_23_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_23_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1
      ^ state_2_42_1_lpi_4 ^ state_0_42_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_51_sva_1
      ^ state_2_51_1_lpi_4;
  assign mux1h_77_nl = MUX1HOT_s_1_5_2(state_xor_121_nl, state_0_23_sva_2_mx0w1,
      state_xor_122_nl, data_out_rsci_idat_23, state_xor_123_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_124_nl = xor_cse_414 ^ xor_cse_909 ^ xor_cse_1009 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_20
      ^ Encrypt_Top_sbox_and_1_cse_52_sva_1 ^ Encrypt_Top_sbox_and_2_cse_52_sva_1;
  assign state_xor_125_nl = xor_cse_915 ^ xor_cse_14 ^ xor_cse_316 ^ Encrypt_Top_sbox_1_and_cse_24_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_24_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1;
  assign state_xor_126_nl = state_0_52_lpi_6 ^ xor_cse_316 ^ xor_cse_920 ^ xor_cse_726
      ^ Encrypt_Top_sbox_1_and_cse_24_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_24_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1 ^ state_0_43_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_52_sva_1
      ^ state_2_52_1_lpi_4;
  assign mux1h_78_nl = MUX1HOT_s_1_5_2(state_xor_124_nl, state_0_24_sva_2_mx0w1,
      state_xor_125_nl, data_out_rsci_idat_24, state_xor_126_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_127_nl = xor_cse_427 ^ xor_cse_923 ^ xor_cse_1016 ^ xor_cse_1017;
  assign state_xor_128_nl = state_0_53_lpi_6 ^ xor_cse_325 ^ xor_cse_29 ^ xor_cse_160
      ^ xor_cse_1018 ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1 ^ state_0_44_lpi_6 ^
      Encrypt_Top_sbox_1_and_1_cse_53_sva_1 ^ state_2_53_1_lpi_4;
  assign state_xor_129_nl = state_0_53_lpi_6 ^ xor_cse_325 ^ xor_cse_1018 ^ xor_cse_568
      ^ xor_cse_734 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1 ^ state_0_44_lpi_6 ^
      Encrypt_Top_sbox_3_and_1_cse_53_sva_1 ^ state_2_53_1_lpi_4;
  assign mux1h_79_nl = MUX1HOT_s_1_5_2(state_xor_127_nl, state_0_25_sva_2_mx0w1,
      state_xor_128_nl, data_out_rsci_idat_25, state_xor_129_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_130_nl = Encrypt_Top_sbox_and_2_cse_54_sva_1 ^ xor_cse_1021 ^
      xor_cse_935 ^ xor_cse_448 ^ Encrypt_Top_sbox_and_1_cse_26_sva_1 ^ state_2_26_1_lpi_4
      ^ state_0_26_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_13 ^ Encrypt_Top_sbox_and_1_cse_45_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_45_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_22
      ^ Encrypt_Top_sbox_and_1_cse_54_sva_1;
  assign state_xor_131_nl = xor_cse_450 ^ xor_cse_43 ^ xor_cse_168 ^ Encrypt_Top_sbox_1_and_1_cse_45_sva_1
      ^ state_2_45_1_lpi_4 ^ state_0_45_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1;
  assign state_xor_132_nl = xor_cse_450 ^ xor_cse_740 ^ xor_cse_944 ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1 ^ state_0_45_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1
      ^ state_2_54_1_lpi_4 ^ state_0_54_lpi_6;
  assign mux1h_80_nl = MUX1HOT_s_1_5_2(state_xor_130_nl, state_0_26_sva_2_mx0w1,
      state_xor_131_nl, data_out_rsci_idat_26, state_xor_132_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_133_nl = xor_cse_947 ^ xor_cse_1030 ^ xor_cse_1031 ^ Encrypt_Top_sbox_and_1_cse_27_sva_1
      ^ state_2_27_1_lpi_4 ^ state_0_27_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_23
      ^ Encrypt_Top_sbox_and_1_cse_55_sva_1 ^ Encrypt_Top_sbox_and_2_cse_55_sva_1;
  assign state_xor_134_nl = xor_cse_1034 ^ xor_cse_57 ^ xor_cse_181 ^ Encrypt_Top_sbox_1_and_1_cse_46_sva_1
      ^ state_2_46_1_lpi_4 ^ state_0_46_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_55_sva_1
      ^ xor_cse_1037;
  assign state_xor_135_nl = xor_cse_1034 ^ xor_cse_746 ^ xor_cse_604 ^ Encrypt_Top_sbox_3_and_1_cse_46_sva_1
      ^ state_2_46_1_lpi_4 ^ state_0_46_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1
      ^ xor_cse_1037;
  assign mux1h_81_nl = MUX1HOT_s_1_5_2(state_xor_133_nl, state_0_27_sva_2_mx0w1,
      state_xor_134_nl, data_out_rsci_idat_27, state_xor_135_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_136_nl = Encrypt_Top_sbox_and_2_cse_56_sva_1 ^ xor_cse_1041 ^
      xor_cse_961 ^ xor_cse_354 ^ Encrypt_Top_sbox_and_1_cse_28_sva_1 ^ state_2_28_1_lpi_4
      ^ state_0_28_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_15 ^ Encrypt_Top_sbox_and_1_cse_47_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_47_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_24
      ^ Encrypt_Top_sbox_and_1_cse_56_sva_1;
  assign state_xor_137_nl = xor_cse_356 ^ xor_cse_73 ^ xor_cse_192 ^ Encrypt_Top_sbox_1_and_1_cse_47_sva_1
      ^ state_2_47_1_lpi_4 ^ state_0_47_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_56_sva_1
      ^ xor_cse_1046;
  assign state_xor_138_nl = xor_cse_356 ^ xor_cse_967 ^ xor_cse_752 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1 ^ state_0_47_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_56_sva_1
      ^ xor_cse_1046;
  assign mux1h_82_nl = MUX1HOT_s_1_5_2(state_xor_136_nl, state_0_28_sva_2_mx0w1,
      state_xor_137_nl, data_out_rsci_idat_28, state_xor_138_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_139_nl = Encrypt_Top_sbox_and_2_cse_57_sva_1 ^ xor_cse_1050 ^
      xor_cse_970 ^ xor_cse_366 ^ Encrypt_Top_sbox_and_1_cse_29_sva_1 ^ state_2_29_1_lpi_4
      ^ state_0_29_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_16 ^ Encrypt_Top_sbox_and_1_cse_48_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_48_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_25
      ^ Encrypt_Top_sbox_and_1_cse_57_sva_1;
  assign state_xor_140_nl = xor_cse_368 ^ xor_cse_85 ^ xor_cse_201 ^ Encrypt_Top_sbox_1_and_1_cse_48_sva_1
      ^ state_2_48_1_lpi_4 ^ state_0_48_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1
      ^ xor_cse_1055;
  assign state_xor_141_nl = xor_cse_368 ^ xor_cse_977 ^ xor_cse_470 ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1 ^ state_0_48_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1
      ^ xor_cse_1055;
  assign mux1h_83_nl = MUX1HOT_s_1_5_2(state_xor_139_nl, state_0_29_sva_2_mx0w1,
      state_xor_140_nl, data_out_rsci_idat_29, state_xor_141_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_142_nl = Encrypt_Top_sbox_and_2_cse_58_sva_1 ^ xor_cse_1059 ^
      xor_cse_981 ^ xor_cse_379 ^ Encrypt_Top_sbox_and_1_cse_30_sva_1 ^ state_2_30_1_lpi_4
      ^ state_0_30_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_17 ^ Encrypt_Top_sbox_and_1_cse_49_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_49_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_26
      ^ Encrypt_Top_sbox_and_1_cse_58_sva_1;
  assign state_xor_143_nl = xor_cse_871 ^ xor_cse_100 ^ xor_cse_214 ^ Encrypt_Top_sbox_1_and_1_cse_49_sva_1
      ^ state_2_49_1_lpi_4 ^ state_0_49_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_58_sva_1
      ^ xor_cse_1064;
  assign state_xor_144_nl = xor_cse_871 ^ xor_cse_480 ^ xor_cse_702 ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1
      ^ state_2_49_1_lpi_4 ^ state_0_49_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1
      ^ xor_cse_1064;
  assign mux1h_84_nl = MUX1HOT_s_1_5_2(state_xor_142_nl, state_0_30_sva_2_mx0w1,
      state_xor_143_nl, data_out_rsci_idat_30, state_xor_144_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_145_nl = Encrypt_Top_sbox_and_2_cse_59_sva_1 ^ xor_cse_1068 ^
      xor_cse_990 ^ xor_cse_390 ^ Encrypt_Top_sbox_and_1_cse_31_sva_1 ^ state_2_31_1_lpi_4
      ^ state_0_31_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_18 ^ Encrypt_Top_sbox_and_1_cse_50_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_50_sva_1 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_27
      ^ Encrypt_Top_sbox_and_1_cse_59_sva_1;
  assign state_xor_146_nl = xor_cse_393 ^ xor_cse_115 ^ xor_cse_224 ^ Encrypt_Top_sbox_1_and_1_cse_50_sva_1
      ^ state_2_50_1_lpi_4 ^ state_0_50_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_59_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1 ^ state_0_59_lpi_6;
  assign state_xor_147_nl = xor_cse_393 ^ xor_cse_996 ^ xor_cse_492 ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_50_sva_1 ^ state_0_50_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1
      ^ state_2_59_1_lpi_4 ^ state_0_59_lpi_6;
  assign mux1h_85_nl = MUX1HOT_s_1_5_2(state_xor_145_nl, state_0_31_sva_2_mx0w1,
      state_xor_146_nl, data_out_rsci_idat_31, state_xor_147_nl, {(fsm_output[1])
      , (fsm_output[3]) , and_24_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_148_nl = xor_cse_1077 ^ xor_cse_400 ^ xor_cse_1000 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_19
      ^ Encrypt_Top_sbox_and_1_cse_51_sva_1 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1;
  assign state_xor_149_nl = xor_cse ^ xor_cse_3 ^ xor_cse_4 ^ xor_cse_5 ^ state_2_32_1_lpi_4
      ^ state_0_32_lpi_6;
  assign state_xor_150_nl = xor_cse_895 ^ xor_cse_499 ^ xor_cse_717 ^ Encrypt_Top_sbox_3_and_1_cse_51_sva_1
      ^ state_2_51_1_lpi_4 ^ state_0_51_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1
      ^ xor_cse_1085;
  assign mux1h_86_nl = MUX1HOT_s_1_6_2(state_xor_148_nl, ADLEN_ADLEN_xor_2_itm_mx0w0,
      state_xor_149_nl, state_0_4_sva_4_mx0w4, state_0_4_lpi_6, state_xor_150_nl,
      {(fsm_output[1]) , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xor_151_nl = xor_cse_1086 ^ xor_cse_1009 ^ xor_cse_419 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_1
      ^ Encrypt_Top_sbox_and_1_cse_33_sva_1 ^ Encrypt_Top_sbox_and_2_cse_33_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_20 ^ Encrypt_Top_sbox_and_1_cse_52_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_52_sva_1;
  assign state_xor_152_nl = xor_cse_14 ^ xor_cse_17 ^ xor_cse_18 ^ xor_cse_19 ^ state_2_33_1_lpi_4
      ^ state_0_33_lpi_6;
  assign state_xor_153_nl = xor_cse_906 ^ xor_cse_515 ^ xor_cse_726 ^ Encrypt_Top_sbox_3_and_1_cse_52_sva_1
      ^ state_2_52_1_lpi_4 ^ state_0_52_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_61_sva_1
      ^ xor_cse_1095;
  assign mux1h_87_nl = MUX1HOT_s_1_6_2(state_xor_151_nl, ADLEN_ADLEN_xor_4_itm_mx0w0,
      state_xor_152_nl, state_0_5_sva_4_mx0w4, state_0_5_lpi_6, state_xor_153_nl,
      {(fsm_output[1]) , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xor_154_nl = xor_cse_1096 ^ xor_cse_1016 ^ xor_cse_431 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_2
      ^ Encrypt_Top_sbox_and_1_cse_34_sva_1 ^ Encrypt_Top_sbox_and_2_cse_34_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_21 ^ Encrypt_Top_sbox_and_1_cse_53_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_53_sva_1;
  assign state_xor_155_nl = Encrypt_Top_sbox_1_and_1_cse_53_sva_1 ^ xor_cse_28 ^
      xor_cse_29 ^ xor_cse_30 ^ xor_cse_31 ^ xor_cse_32;
  assign state_xor_156_nl = state_0_62_lpi_6 ^ xor_cse_439 ^ xor_cse_521 ^ xor_cse_734
      ^ xor_cse_32 ^ Encrypt_Top_sbox_3_and_1_cse_34_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_53_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1 ^ state_2_62_1_lpi_4;
  assign mux1h_88_nl = MUX1HOT_s_1_6_2(state_xor_154_nl, ADLEN_ADLEN_xor_6_itm_mx0w0,
      state_xor_155_nl, state_0_6_sva_4_mx0w4, state_0_6_lpi_6, state_xor_156_nl,
      {(fsm_output[1]) , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xor_157_nl = xor_cse_445 ^ xor_cse_1103 ^ xor_cse_1021 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_22
      ^ Encrypt_Top_sbox_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_and_2_cse_54_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_31 ^ Encrypt_Top_sbox_and_1_cse_63_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_63_sva_1;
  assign state_xor_158_nl = xor_cse_46 ^ xor_cse_47 ^ xor_cse_41 ^ xor_cse_43;
  assign state_xor_159_nl = xor_cse_457 ^ xor_cse_740 ^ xor_cse_527 ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1
      ^ state_2_54_1_lpi_4 ^ state_0_54_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1
      ^ xor_cse_1108;
  assign mux1h_89_nl = MUX1HOT_s_1_6_2(state_xor_157_nl, ADLEN_ADLEN_xor_8_itm_mx0w0,
      state_xor_158_nl, state_0_7_sva_4_mx0w4, state_0_7_lpi_6, state_xor_159_nl,
      {(fsm_output[1]) , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xor_160_nl = xor_cse_351 ^ xor_cse_1030 ^ xor_cse_936 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_4
      ^ Encrypt_Top_sbox_and_1_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_36_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_23 ^ Encrypt_Top_sbox_and_1_cse_55_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_55_sva_1 ^ plaintext_31_0_sva_0;
  assign state_xor_161_nl = xor_cse_59 ^ xor_cse_61 ^ xor_cse_55 ^ xor_cse_359;
  assign state_xor_162_nl = xor_cse_59 ^ xor_cse_60 ^ xor_cse_61 ^ xor_cse_55;
  assign state_xor_164_nl = xor_cse_56 ^ xor_cse_943 ^ xor_cse_746 ^ xor_cse_360
      ^ Encrypt_Top_sbox_3_and_1_cse_36_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1
      ^ state_0_36_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1 ^ xor_cse_1037;
  assign mux1h_90_nl = MUX1HOT_s_1_7_2(state_xor_160_nl, ADLEN_ADLEN_xor_10_itm_mx0w0,
      state_xor_161_nl, state_xor_162_nl, state_0_8_sva_3_mx0w5, state_0_8_lpi_6,
      state_xor_164_nl, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse
      , and_90_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_165_nl = xor_cse_363 ^ xor_cse_1041 ^ xor_cse_950 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_5
      ^ Encrypt_Top_sbox_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_and_2_cse_37_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_24 ^ Encrypt_Top_sbox_and_1_cse_56_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_56_sva_1 ^ plaintext_31_0_sva_1;
  assign state_xor_166_nl = xor_cse_70 ^ xor_cse_73 ^ xor_cse_74 ^ xor_cse_75 ^ state_2_37_1_lpi_4
      ^ state_0_37_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_1_sva_1 ^ state_2_1_1_lpi_4
      ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]) ^ state_0_1_lpi_6;
  assign state_xor_167_nl = xor_cse_73 ^ xor_cse_74 ^ xor_cse_75 ^ xor_cse_69;
  assign state_xor_169_nl = xor_cse_70 ^ xor_cse_958 ^ xor_cse_752 ^ xor_cse_373
      ^ Encrypt_Top_sbox_3_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1
      ^ state_0_37_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_56_sva_1 ^ xor_cse_1046;
  assign mux1h_91_nl = MUX1HOT_s_1_7_2(state_xor_165_nl, ADLEN_ADLEN_xor_12_itm_mx0w0,
      state_xor_166_nl, state_xor_167_nl, state_0_9_sva_3_mx0w5, state_0_9_lpi_6,
      state_xor_169_nl, {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse
      , and_90_cse , (fsm_output[13]) , (fsm_output[14])});
  assign state_xor_170_nl = xor_cse_858 ^ xor_cse_376 ^ xor_cse_1050 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_25
      ^ Encrypt_Top_sbox_and_1_cse_57_sva_1 ^ Encrypt_Top_sbox_and_2_cse_57_sva_1
      ^ plaintext_31_0_sva_2;
  assign state_xor_171_nl = xor_cse_87 ^ xor_cse_89 ^ xor_cse_382 ^ xor_cse_83;
  assign state_xor_172_nl = xor_cse_87 ^ xor_cse_88 ^ xor_cse_89 ^ xor_cse_83;
  assign state_xor_173_nl = xor_cse_866 ^ xor_cse_84 ^ xor_cse_470 ^ xor_cse_385
      ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1 ^ state_2_57_1_lpi_4 ^ state_0_57_lpi_6;
  assign mux1h_92_nl = MUX1HOT_s_1_6_2(state_xor_170_nl, ADLEN_ADLEN_xor_14_itm_mx0w0,
      state_xor_171_nl, state_xor_172_nl, ciphertext_38_sva_mx0w2, state_xor_173_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_174_nl = xor_cse_389 ^ xor_cse_1059 ^ xor_cse_867 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_7
      ^ Encrypt_Top_sbox_and_1_cse_39_sva_1 ^ Encrypt_Top_sbox_and_2_cse_39_sva_1
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_26 ^ Encrypt_Top_sbox_and_1_cse_58_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_58_sva_1 ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_3
      ^ Encrypt_Top_sbox_and_1_cse_3_sva_1 ^ Encrypt_Top_sbox_and_2_cse_3_sva_1 ^
      plaintext_31_0_sva_3;
  assign state_xor_175_nl = xor_cse_97 ^ xor_cse_1134 ^ xor_cse_100 ^ Encrypt_Top_sbox_1_and_1_cse_3_sva_1
      ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3]);
  assign state_xor_176_nl = xor_cse_102 ^ xor_cse_103 ^ xor_cse_97 ^ xor_cse_99;
  assign state_xor_177_nl = xor_cse_1134 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3])
      ^ xor_cse_480 ^ xor_cse_875 ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_39_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_3_sva_1;
  assign mux1h_93_nl = MUX1HOT_s_1_6_2(state_xor_174_nl, ADLEN_ADLEN_xor_16_itm_mx0w0,
      state_xor_175_nl, state_xor_176_nl, ciphertext_39_sva_mx0w2, state_xor_177_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_178_nl = xor_cse_877 ^ xor_cse_405 ^ xor_cse_1068 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_27
      ^ Encrypt_Top_sbox_and_1_cse_59_sva_1 ^ Encrypt_Top_sbox_and_2_cse_59_sva_1
      ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_4 ^ Encrypt_Top_sbox_and_1_cse_4_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_4_sva_1 ^ plaintext_31_0_sva_4;
  assign state_xor_179_nl = xor_cse_110 ^ xor_cse_115 ^ xor_cse_113 ^ xor_cse_1144
      ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1
      ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign state_xor_180_nl = xor_cse_115 ^ xor_cse_116 ^ xor_cse_110 ^ xor_cse_112;
  assign state_xor_181_nl = xor_cse_111 ^ xor_cse_492 ^ xor_cse_635 ^ xor_cse_1144
      ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1
      ^ state_2_59_1_lpi_4 ^ state_0_59_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_4_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4]);
  assign mux1h_94_nl = MUX1HOT_s_1_6_2(state_xor_178_nl, ADLEN_ADLEN_xor_18_itm_mx0w0,
      state_xor_179_nl, state_xor_180_nl, ciphertext_40_sva_mx0w2, state_xor_181_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_182_nl = plaintext_31_0_sva_5 ^ xor_cse_1077 ^ xor_cse_887 ^ xor_cse_416;
  assign state_xor_183_nl = xor_cse_3 ^ xor_cse_124 ^ xor_cse_127 ^ xor_cse_128 ^
      Encrypt_Top_sbox_2_and_2_cse_41_sva_1 ^ state_0_41_lpi_6 ^ Encrypt_Top_sbox_1_and_1_cse_5_sva_1
      ^ state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5])
      ^ state_0_5_lpi_6;
  assign state_xor_184_nl = xor_cse_3 ^ xor_cse_127 ^ xor_cse_128 ^ xor_cse_123;
  assign state_xor_185_nl = xor_cse_124 ^ xor_cse_897 ^ xor_cse_499 ^ xor_cse_426
      ^ Encrypt_Top_sbox_3_and_1_cse_41_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_41_sva_1
      ^ state_0_41_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1 ^ xor_cse_1085;
  assign mux1h_95_nl = MUX1HOT_s_1_6_2(state_xor_182_nl, ADLEN_ADLEN_xor_20_itm_mx0w0,
      state_xor_183_nl, state_xor_184_nl, ciphertext_41_sva_mx0w2, state_xor_185_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_186_nl = xor_cse_1086 ^ xor_cse_430 ^ xor_cse_899 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_10
      ^ Encrypt_Top_sbox_and_1_cse_42_sva_1 ^ Encrypt_Top_sbox_and_2_cse_42_sva_1
      ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_6 ^ Encrypt_Top_sbox_and_1_cse_6_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_6_sva_1 ^ plaintext_31_0_sva_6;
  assign state_xor_187_nl = xor_cse_17 ^ xor_cse_136 ^ xor_cse_139 ^ xor_cse_140
      ^ xor_cse_435 ^ xor_cse_905;
  assign state_xor_188_nl = xor_cse_17 ^ xor_cse_139 ^ xor_cse_140 ^ xor_cse_135;
  assign state_xor_189_nl = xor_cse_136 ^ xor_cse_515 ^ xor_cse_651 ^ xor_cse_441
      ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1 ^ state_2_42_1_lpi_4 ^ state_0_42_lpi_6
      ^ Encrypt_Top_sbox_3_and_1_cse_61_sva_1 ^ xor_cse_1095;
  assign mux1h_96_nl = MUX1HOT_s_1_6_2(state_xor_186_nl, ADLEN_ADLEN_xor_22_itm_mx0w0,
      state_xor_187_nl, state_xor_188_nl, ciphertext_42_sva_mx0w2, state_xor_189_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_190_nl = plaintext_31_0_sva_7 ^ xor_cse_1096 ^ xor_cse_443 ^ xor_cse_909;
  assign state_xor_191_nl = xor_cse_148 ^ xor_cse_28 ^ xor_cse_151 ^ xor_cse_152
      ^ xor_cse_452 ^ state_2_43_1_lpi_4 ^ state_0_43_lpi_6;
  assign state_xor_192_nl = xor_cse_28 ^ xor_cse_151 ^ xor_cse_152 ^ xor_cse_147;
  assign state_xor_193_nl = xor_cse_148 ^ xor_cse_920 ^ xor_cse_521 ^ xor_cse_456
      ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_43_sva_1
      ^ state_0_43_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1 ^ state_2_62_1_lpi_4
      ^ state_0_62_lpi_6;
  assign mux1h_97_nl = MUX1HOT_s_1_6_2(state_xor_190_nl, ADLEN_ADLEN_xor_24_itm_mx0w0,
      state_xor_191_nl, state_xor_192_nl, ciphertext_43_sva_mx0w2, state_xor_193_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_197_nl = xor_cse_1171 ^ xor_cse_351 ^ xor_cse_935 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_13
      ^ Encrypt_Top_sbox_and_1_cse_45_sva_1 ^ Encrypt_Top_sbox_and_2_cse_45_sva_1
      ^ plaintext_31_0_sva_0;
  assign state_xor_198_nl = xor_cse_170 ^ xor_cse_171 ^ xor_cse_359 ^ xor_cse_167;
  assign state_xor_199_nl = xor_cse_170 ^ xor_cse_60 ^ xor_cse_171 ^ xor_cse_167;
  assign state_xor_200_nl = xor_cse_56 ^ xor_cse_506 ^ xor_cse_944 ^ xor_cse_360
      ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_45_sva_1
      ^ state_0_45_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_9_sva_1 ^ state_2_9_1_lpi_4
      ^ state_0_9_lpi_6;
  assign mux1h_99_nl = MUX1HOT_s_1_6_2(state_xor_197_nl, ADLEN_ADLEN_xor_28_itm_mx0w0,
      state_xor_198_nl, state_xor_199_nl, ciphertext_45_sva_mx0w2, state_xor_200_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_201_nl = xor_cse_947 ^ xor_cse_363 ^ xor_cse_861 ^ plaintext_31_0_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_10_sva_1 ^ state_2_10_1_lpi_4 ^ state_0_10_lpi_6;
  assign state_xor_202_nl = xor_cse_177 ^ state_0_1_lpi_6 ^ xor_cse_181 ^ Encrypt_Top_sbox_1_and_1_cse_46_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_1_sva_1 ^ state_2_1_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1]);
  assign state_xor_203_nl = Encrypt_Top_sbox_1_and_1_cse_46_sva_1 ^ xor_cse_181 ^
      xor_cse_71 ^ xor_cse_177;
  assign state_xor_204_nl = Encrypt_Top_sbox_3_and_1_cse_46_sva_1 ^ xor_cse_604 ^
      xor_cse_373 ^ xor_cse_177;
  assign mux1h_100_nl = MUX1HOT_s_1_6_2(state_xor_201_nl, ADLEN_ADLEN_xor_30_itm_mx0w0,
      state_xor_202_nl, state_xor_203_nl, ciphertext_46_sva_mx0w2, state_xor_204_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_205_nl = xor_cse_376 ^ xor_cse_961 ^ xor_cse_868 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_15
      ^ Encrypt_Top_sbox_and_1_cse_47_sva_1 ^ Encrypt_Top_sbox_and_2_cse_47_sva_1
      ^ plaintext_31_0_sva_2 ^ Encrypt_Top_sbox_and_1_cse_11_sva_1 ^ state_2_11_1_lpi_4
      ^ state_0_11_lpi_6;
  assign state_xor_206_nl = state_2_47_1_lpi_4 ^ xor_cse_192 ^ xor_cse_382 ^ xor_cse_188;
  assign state_xor_207_nl = state_2_47_1_lpi_4 ^ xor_cse_192 ^ xor_cse_88 ^ xor_cse_188;
  assign state_xor_208_nl = xor_cse_190 ^ xor_cse_189 ^ xor_cse_84 ^ xor_cse_967
      ^ xor_cse_385 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_47_sva_1;
  assign mux1h_101_nl = MUX1HOT_s_1_6_2(state_xor_205_nl, ADLEN_ADLEN_xor_32_itm_mx0w0,
      state_xor_206_nl, state_xor_207_nl, ciphertext_47_sva_mx0w2, state_xor_208_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_209_nl = xor_cse_389 ^ xor_cse_970 ^ xor_cse_880 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_16
      ^ Encrypt_Top_sbox_and_1_cse_48_sva_1 ^ Encrypt_Top_sbox_and_2_cse_48_sva_1
      ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_3 ^ Encrypt_Top_sbox_and_1_cse_3_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_3_sva_1 ^ plaintext_31_0_sva_3 ^ Encrypt_Top_sbox_and_1_cse_12_sva_1
      ^ xor_cse_1187;
  assign state_xor_210_nl = Encrypt_Top_sbox_1_and_1_cse_3_sva_1 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3])
      ^ xor_cse_1188 ^ xor_cse_200;
  assign state_xor_211_nl = xor_cse_204 ^ xor_cse_102 ^ xor_cse_103 ^ xor_cse_200;
  assign state_xor_212_nl = xor_cse_1188 ^ xor_cse_202 ^ xor_cse_977 ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_48_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_3_sva_1
      ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[3]);
  assign mux1h_102_nl = MUX1HOT_s_1_6_2(state_xor_209_nl, ADLEN_ADLEN_xor_34_itm_mx0w0,
      state_xor_210_nl, state_xor_211_nl, ciphertext_48_sva_mx0w2, state_xor_212_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_213_nl = xor_cse_405 ^ xor_cse_981 ^ xor_cse_890 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_17
      ^ Encrypt_Top_sbox_and_1_cse_49_sva_1 ^ Encrypt_Top_sbox_and_2_cse_49_sva_1
      ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_4 ^ Encrypt_Top_sbox_and_1_cse_4_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_4_sva_1 ^ plaintext_31_0_sva_4 ^ Encrypt_Top_sbox_and_1_cse_13_sva_1
      ^ xor_cse_1193;
  assign state_xor_214_nl = xor_cse_210 ^ state_0_4_lpi_6 ^ xor_cse_214 ^ Encrypt_Top_sbox_1_and_1_cse_49_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1 ^ state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4]);
  assign state_xor_215_nl = Encrypt_Top_sbox_1_and_1_cse_49_sva_1 ^ xor_cse_214 ^
      xor_cse_116 ^ xor_cse_210;
  assign state_xor_216_nl = xor_cse_210 ^ state_0_4_lpi_6 ^ xor_cse_702 ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_4_sva_1 ^ state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[4]);
  assign mux1h_103_nl = MUX1HOT_s_1_6_2(state_xor_213_nl, ADLEN_ADLEN_xor_36_itm_mx0w0,
      state_xor_214_nl, state_xor_215_nl, ciphertext_49_sva_mx0w2, state_xor_216_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_217_nl = xor_cse_416 ^ xor_cse_990 ^ xor_cse_900 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_18
      ^ Encrypt_Top_sbox_and_1_cse_50_sva_1 ^ Encrypt_Top_sbox_and_2_cse_50_sva_1
      ^ plaintext_31_0_sva_5 ^ Encrypt_Top_sbox_and_1_cse_14_sva_1 ^ state_2_14_1_lpi_4
      ^ state_0_14_lpi_6;
  assign state_xor_218_nl = xor_cse_220 ^ state_0_5_lpi_6 ^ xor_cse_224 ^ state_2_50_1_lpi_4
      ^ Encrypt_Top_sbox_1_and_1_cse_5_sva_1 ^ state_2_5_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]);
  assign state_xor_219_nl = state_2_50_1_lpi_4 ^ xor_cse_224 ^ xor_cse_125 ^ xor_cse_220;
  assign state_xor_220_nl = xor_cse_222 ^ xor_cse_221 ^ xor_cse_124 ^ xor_cse_996
      ^ xor_cse_426 ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1 ^ Encrypt_Top_sbox_3_and_2_cse_50_sva_1;
  assign mux1h_104_nl = MUX1HOT_s_1_6_2(state_xor_217_nl, ADLEN_ADLEN_xor_38_itm_mx0w0,
      state_xor_218_nl, state_xor_219_nl, ciphertext_50_sva_mx0w2, state_xor_220_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_221_nl = xor_cse_430 ^ xor_cse_1000 ^ xor_cse_912 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_19
      ^ Encrypt_Top_sbox_and_1_cse_51_sva_1 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1
      ^ Encrypt_Top_sbox_and_cse_31_0_sva_1_6 ^ Encrypt_Top_sbox_and_1_cse_6_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_6_sva_1 ^ plaintext_31_0_sva_6 ^ Encrypt_Top_sbox_and_1_cse_15_sva_1
      ^ state_2_15_1_lpi_4 ^ state_0_15_lpi_6;
  assign state_xor_222_nl = Encrypt_Top_sbox_1_and_1_cse_51_sva_1 ^ xor_cse_1 ^ xor_cse_230
      ^ xor_cse_435;
  assign state_xor_223_nl = Encrypt_Top_sbox_1_and_1_cse_51_sva_1 ^ xor_cse_1 ^ xor_cse_137
      ^ xor_cse_230;
  assign state_xor_224_nl = Encrypt_Top_sbox_3_and_1_cse_51_sva_1 ^ xor_cse_717 ^
      xor_cse_441 ^ xor_cse_230;
  assign mux1h_105_nl = MUX1HOT_s_1_6_2(state_xor_221_nl, ADLEN_ADLEN_xor_40_itm_mx0w0,
      state_xor_222_nl, state_xor_223_nl, ciphertext_51_sva_mx0w2, state_xor_224_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_225_nl = xor_cse_443 ^ xor_cse_1009 ^ xor_cse_926 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_20
      ^ Encrypt_Top_sbox_and_1_cse_52_sva_1 ^ Encrypt_Top_sbox_and_2_cse_52_sva_1
      ^ plaintext_31_0_sva_7 ^ xor_cse_927;
  assign state_xor_226_nl = Encrypt_Top_sbox_1_and_1_cse_52_sva_1 ^ xor_cse_15 ^
      xor_cse_241 ^ xor_cse_452;
  assign state_xor_227_nl = Encrypt_Top_sbox_1_and_1_cse_52_sva_1 ^ xor_cse_15 ^
      xor_cse_149 ^ xor_cse_241;
  assign state_xor_228_nl = Encrypt_Top_sbox_3_and_1_cse_52_sva_1 ^ xor_cse_726 ^
      xor_cse_456 ^ xor_cse_241;
  assign mux1h_106_nl = MUX1HOT_s_1_6_2(state_xor_225_nl, ADLEN_ADLEN_xor_42_itm_mx0w0,
      state_xor_226_nl, state_xor_227_nl, ciphertext_52_sva_mx0w2, state_xor_228_nl,
      {(fsm_output[1]) , (fsm_output[2]) , (fsm_output[4]) , and_21_cse , and_90_cse
      , (fsm_output[14])});
  assign state_xor_194_nl = xor_cse_1161 ^ xor_cse_923 ^ xor_cse_1103 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_31
      ^ Encrypt_Top_sbox_and_1_cse_63_sva_1 ^ Encrypt_Top_sbox_and_2_cse_63_sva_1;
  assign state_xor_195_nl = xor_cse_41 ^ xor_cse_159 ^ xor_cse_160 ^ xor_cse_161
      ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1 ^ state_0_44_lpi_6;
  assign state_xor_196_nl = xor_cse_1167 ^ xor_cse_527 ^ xor_cse_568 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1
      ^ state_2_44_1_lpi_4 ^ state_0_44_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1
      ^ xor_cse_1108;
  assign mux1h_98_nl = MUX1HOT_s_1_5_2(state_xor_194_nl, ADLEN_ADLEN_xor_26_itm_mx0w0,
      state_xor_195_nl, ciphertext_44_sva_mx0w2, state_xor_196_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_229_nl = xor_cse_932 ^ xor_cse_1161 ^ xor_cse_1016 ^ xor_cse_1017;
  assign state_xor_230_nl = xor_cse_251 ^ xor_cse_29 ^ xor_cse_159 ^ xor_cse_254
      ^ state_2_8_1_lpi_4 ^ state_0_8_lpi_6;
  assign state_xor_231_nl = xor_cse_251 ^ xor_cse_1167 ^ xor_cse_734 ^ Encrypt_Top_sbox_3_and_1_cse_53_sva_1
      ^ state_2_53_1_lpi_4 ^ state_0_53_lpi_6;
  assign mux1h_107_nl = MUX1HOT_s_1_5_2(state_xor_229_nl, ADLEN_ADLEN_xor_44_itm_mx0w0,
      state_xor_230_nl, ciphertext_53_sva_mx0w2, state_xor_231_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_232_nl = xor_cse_1171 ^ xor_cse_1021 ^ xor_cse_951 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_22
      ^ Encrypt_Top_sbox_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_and_2_cse_54_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_18_sva_1 ^ state_2_18_1_lpi_4 ^ state_0_18_lpi_6;
  assign state_xor_233_nl = xor_cse_262 ^ xor_cse_44 ^ xor_cse_170 ^ xor_cse_265
      ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_9_sva_1;
  assign state_xor_234_nl = xor_cse_262 ^ xor_cse_740 ^ xor_cse_506 ^ xor_cse_265
      ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_9_sva_1;
  assign mux1h_108_nl = MUX1HOT_s_1_5_2(state_xor_232_nl, ADLEN_ADLEN_xor_46_itm_mx0w0,
      state_xor_233_nl, ciphertext_54_sva_mx0w2, state_xor_234_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_235_nl = xor_cse_349 ^ xor_cse_1030 ^ xor_cse_861 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_23
      ^ Encrypt_Top_sbox_and_1_cse_55_sva_1 ^ Encrypt_Top_sbox_and_2_cse_55_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_10_sva_1 ^ state_2_10_1_lpi_4 ^ state_0_10_lpi_6;
  assign state_xor_236_nl = xor_cse_272 ^ xor_cse_274 ^ xor_cse_57 ^ xor_cse_275
      ^ Encrypt_Top_sbox_1_and_1_cse_55_sva_1 ^ state_0_55_lpi_6;
  assign state_xor_237_nl = xor_cse_272 ^ xor_cse_274 ^ xor_cse_746 ^ xor_cse_275
      ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1 ^ state_0_55_lpi_6;
  assign mux1h_109_nl = MUX1HOT_s_1_5_2(state_xor_235_nl, ADLEN_ADLEN_xor_48_itm_mx0w0,
      state_xor_236_nl, ciphertext_55_sva_mx0w2, state_xor_237_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_238_nl = xor_cse_361 ^ xor_cse_1041 ^ xor_cse_868 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_24
      ^ Encrypt_Top_sbox_and_1_cse_56_sva_1 ^ Encrypt_Top_sbox_and_2_cse_56_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_11_sva_1 ^ state_2_11_1_lpi_4 ^ state_0_11_lpi_6;
  assign state_xor_239_nl = xor_cse_280 ^ xor_cse_282 ^ xor_cse_73 ^ xor_cse_283
      ^ Encrypt_Top_sbox_1_and_1_cse_56_sva_1 ^ state_0_56_lpi_6;
  assign state_xor_240_nl = xor_cse_280 ^ xor_cse_282 ^ xor_cse_752 ^ xor_cse_283
      ^ Encrypt_Top_sbox_3_and_1_cse_56_sva_1 ^ state_0_56_lpi_6;
  assign mux1h_110_nl = MUX1HOT_s_1_5_2(state_xor_238_nl, ADLEN_ADLEN_xor_50_itm_mx0w0,
      state_xor_239_nl, ciphertext_56_sva_mx0w2, state_xor_240_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_241_nl = xor_cse_374 ^ xor_cse_1050 ^ xor_cse_880 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_25
      ^ Encrypt_Top_sbox_and_1_cse_57_sva_1 ^ Encrypt_Top_sbox_and_2_cse_57_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_12_sva_1 ^ xor_cse_1187;
  assign state_xor_242_nl = xor_cse_288 ^ xor_cse_290 ^ xor_cse_85 ^ xor_cse_291
      ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1 ^ state_0_57_lpi_6;
  assign state_xor_243_nl = xor_cse_288 ^ xor_cse_290 ^ xor_cse_470 ^ xor_cse_291
      ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1 ^ state_0_57_lpi_6;
  assign mux1h_111_nl = MUX1HOT_s_1_5_2(state_xor_241_nl, ADLEN_ADLEN_xor_52_itm_mx0w0,
      state_xor_242_nl, ciphertext_57_sva_mx0w2, state_xor_243_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_244_nl = xor_cse_386 ^ xor_cse_1059 ^ xor_cse_890 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_26
      ^ Encrypt_Top_sbox_and_1_cse_58_sva_1 ^ Encrypt_Top_sbox_and_2_cse_58_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_13_sva_1 ^ xor_cse_1193;
  assign state_xor_245_nl = xor_cse_297 ^ xor_cse_299 ^ xor_cse_100 ^ xor_cse_300
      ^ Encrypt_Top_sbox_1_and_1_cse_58_sva_1 ^ state_0_58_lpi_6;
  assign state_xor_246_nl = xor_cse_297 ^ xor_cse_299 ^ xor_cse_480 ^ xor_cse_300
      ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1 ^ state_0_58_lpi_6;
  assign mux1h_112_nl = MUX1HOT_s_1_5_2(state_xor_244_nl, ADLEN_ADLEN_xor_54_itm_mx0w0,
      state_xor_245_nl, ciphertext_58_sva_mx0w2, state_xor_246_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_247_nl = xor_cse_402 ^ xor_cse_1068 ^ xor_cse_900 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_27
      ^ Encrypt_Top_sbox_and_1_cse_59_sva_1 ^ Encrypt_Top_sbox_and_2_cse_59_sva_1
      ^ Encrypt_Top_sbox_and_1_cse_14_sva_1 ^ state_2_14_1_lpi_4 ^ state_0_14_lpi_6;
  assign state_xor_248_nl = xor_cse_306 ^ xor_cse_308 ^ xor_cse_115 ^ xor_cse_309
      ^ Encrypt_Top_sbox_1_and_1_cse_59_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1;
  assign state_xor_249_nl = xor_cse_306 ^ xor_cse_308 ^ xor_cse_492 ^ xor_cse_309
      ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1 ^ state_2_59_1_lpi_4;
  assign mux1h_113_nl = MUX1HOT_s_1_5_2(state_xor_247_nl, ADLEN_ADLEN_xor_56_itm_mx0w0,
      state_xor_248_nl, ciphertext_59_sva_mx0w2, state_xor_249_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_250_nl = xor_cse_1077 ^ xor_cse_414 ^ xor_cse_912 ^ Encrypt_Top_sbox_and_1_cse_15_sva_1
      ^ state_2_15_1_lpi_4 ^ state_0_15_lpi_6;
  assign state_xor_251_nl = xor_cse_315 ^ xor_cse_3 ^ xor_cse_318 ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_60_sva_1 ^ state_1_1_63_32_lpi_4_28;
  assign state_xor_252_nl = xor_cse_315 ^ xor_cse_499 ^ xor_cse_318 ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1
      ^ state_2_60_1_lpi_4 ^ state_0_60_lpi_6;
  assign mux1h_114_nl = MUX1HOT_s_1_5_2(state_xor_250_nl, ADLEN_ADLEN_xor_58_itm_mx0w0,
      state_xor_251_nl, ciphertext_60_sva_mx0w2, state_xor_252_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_253_nl = xor_cse_1086 ^ xor_cse_427 ^ xor_cse_926 ^ xor_cse_927;
  assign state_xor_254_nl = xor_cse_324 ^ xor_cse_17 ^ xor_cse_327 ^ Encrypt_Top_sbox_1_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_61_sva_1 ^ state_1_1_63_32_lpi_4_29;
  assign state_xor_255_nl = xor_cse_324 ^ xor_cse_515 ^ xor_cse_327 ^ Encrypt_Top_sbox_3_and_1_cse_61_sva_1
      ^ state_2_61_1_lpi_4 ^ state_0_61_lpi_6;
  assign mux1h_115_nl = MUX1HOT_s_1_5_2(state_xor_253_nl, ADLEN_ADLEN_xor_60_itm_mx0w0,
      state_xor_254_nl, ciphertext_61_sva_mx0w2, state_xor_255_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_256_nl = xor_cse_1096 ^ xor_cse_932 ^ xor_cse_448 ^ Encrypt_Top_sbox_and_1_cse_26_sva_1
      ^ state_2_26_1_lpi_4 ^ state_0_26_lpi_6;
  assign state_xor_257_nl = xor_cse_333 ^ xor_cse_28 ^ xor_cse_336 ^ Encrypt_Top_sbox_1_and_1_cse_62_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_62_sva_1 ^ state_1_1_63_32_lpi_4_30;
  assign state_xor_258_nl = xor_cse_333 ^ xor_cse_521 ^ xor_cse_336 ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1
      ^ state_2_62_1_lpi_4 ^ state_0_62_lpi_6;
  assign mux1h_116_nl = MUX1HOT_s_1_5_2(state_xor_256_nl, ADLEN_ADLEN_xor_62_itm_mx0w0,
      state_xor_257_nl, ciphertext_62_sva_mx0w2, state_xor_258_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_259_nl = state_0_27_lpi_6 ^ xor_cse_1103 ^ xor_cse_951 ^ xor_cse_1031
      ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_31 ^ Encrypt_Top_sbox_and_1_cse_63_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_63_sva_1 ^ Encrypt_Top_sbox_and_1_cse_18_sva_1
      ^ state_2_18_1_lpi_4 ^ state_0_18_lpi_6 ^ Encrypt_Top_sbox_and_1_cse_27_sva_1
      ^ state_2_27_1_lpi_4;
  assign state_xor_260_nl = xor_cse_341 ^ xor_cse_343 ^ xor_cse_42 ^ xor_cse_344
      ^ Encrypt_Top_sbox_1_and_1_cse_63_sva_1 ^ state_0_63_lpi_6;
  assign state_xor_261_nl = xor_cse_341 ^ xor_cse_343 ^ xor_cse_527 ^ xor_cse_344
      ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1 ^ state_0_63_lpi_6;
  assign mux1h_117_nl = MUX1HOT_s_1_5_2(state_xor_259_nl, ADLEN_ADLEN_xor_64_itm_mx0w0,
      state_xor_260_nl, ciphertext_63_sva_mx0w2, state_xor_261_nl, {(fsm_output[1])
      , (fsm_output[2]) , or_tmp_913 , and_90_cse , (fsm_output[14])});
  assign state_xor_262_nl = xor_cse_1161 ^ xor_cse_936 ^ xor_cse_1031 ^ Encrypt_Top_sbox_and_1_cse_27_sva_1
      ^ state_2_27_1_lpi_4 ^ state_0_27_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_4
      ^ Encrypt_Top_sbox_and_1_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_36_sva_1;
  assign state_xor_263_nl = xor_cse_1034 ^ xor_cse_1167 ^ xor_cse_943 ^ Encrypt_Top_sbox_3_and_1_cse_36_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_36_sva_1 ^ state_0_36_lpi_6;
  assign mux1h_118_nl = MUX1HOT_s_1_6_2(state_xor_262_nl, state_0_8_sva_2_mx0w1,
      state_0_8_sva_3_mx0w5, ciphertext_36_sva_mx0w2, data_out_rsci_idat_8, state_xor_263_nl,
      {(fsm_output[1]) , (fsm_output[3]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xor_264_nl = xor_cse_1171 ^ xor_cse_950 ^ xor_cse_354 ^ Encrypt_Top_sbox_and_1_cse_28_sva_1
      ^ state_2_28_1_lpi_4 ^ state_0_28_lpi_6 ^ Encrypt_Top_sbox_and_cse_63_32_sva_1_5
      ^ xor_cse_953;
  assign state_xor_265_nl = xor_cse_356 ^ xor_cse_958 ^ xor_cse_506 ^ Encrypt_Top_sbox_3_and_1_cse_9_sva_1
      ^ state_2_9_1_lpi_4 ^ state_0_9_lpi_6 ^ Encrypt_Top_sbox_3_and_1_cse_37_sva_1
      ^ Encrypt_Top_sbox_3_and_2_cse_37_sva_1 ^ state_0_37_lpi_6;
  assign mux1h_119_nl = MUX1HOT_s_1_6_2(state_xor_264_nl, state_0_9_sva_2_mx0w1,
      state_0_9_sva_3_mx0w5, ciphertext_37_sva_mx0w2, data_out_rsci_idat_9, state_xor_265_nl,
      {(fsm_output[1]) , (fsm_output[3]) , or_tmp_913 , and_90_cse , (fsm_output[13])
      , (fsm_output[14])});
  assign state_xnor_152_nl = ~(xor_cse_802 ^ xor_cse_809 ^ xor_cse_1293 ^ plaintext_31_0_sva_0
      ^ plaintext_31_0_sva_1 ^ plaintext_31_0_sva_6);
  assign state_xnor_153_nl = ~(xor_cse_814 ^ xor_cse_808 ^ state_1_1_31_0_lpi_4_0
      ^ state_1_1_31_0_lpi_4_1 ^ Encrypt_Top_sbox_1_and_768 ^ state_4_4_6_lpi_3 ^
      state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6]) ^
      state_1_1_31_0_lpi_4_6);
  assign state_xnor_155_nl = ~(xor_cse_809 ^ xor_cse_817 ^ xor_cse_1303 ^ plaintext_31_0_sva_1
      ^ plaintext_31_0_sva_2 ^ plaintext_31_0_sva_7);
  assign state_xnor_156_nl = ~(xor_cse_814 ^ xor_cse_1306 ^ state_1_1_31_0_lpi_4_1
      ^ Encrypt_Top_sbox_1_and_760 ^ state_4_4_2_lpi_3 ^ state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ state_1_1_31_0_lpi_4_2 ^ state_1_1_31_0_lpi_4_7);
  assign state_xnor_158_nl = ~(xor_cse_817 ^ xor_cse_822 ^ xor_cse_845 ^ plaintext_31_0_sva_2
      ^ plaintext_31_0_sva_3);
  assign xor_69_nl = state_2_2_1_lpi_6 ^ (key4[2]);
  assign state_xnor_159_nl = ~(xor_cse_827 ^ Encrypt_Top_sbox_1_and_760 ^ state_4_4_2_lpi_3
      ^ state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[2])
      ^ state_1_1_31_0_lpi_4_2 ^ state_1_1_31_0_lpi_4_3 ^ Encrypt_Top_sbox_1_and_880
      ^ state_4_4_8_lpi_3 ^ state_2_8_1_lpi_4 ^ state_1_1_63_32_lpi_4_8);
  assign state_xnor_161_nl = ~(xor_cse_822 ^ xor_cse_829 ^ xor_cse_847 ^ plaintext_31_0_sva_3
      ^ plaintext_31_0_sva_4);
  assign xor_67_nl = state_2_3_1_lpi_6 ^ (key4[3]);
  assign state_xnor_162_nl = ~(xor_cse_852 ^ xor_cse_834 ^ xor_cse_827 ^ state_1_1_31_0_lpi_4_3
      ^ state_1_1_31_0_lpi_4_4);
  assign state_xnor_164_nl = ~(xor_cse_829 ^ xor_cse_835 ^ plaintext_31_0_sva_4 ^
      plaintext_31_0_sva_5 ^ xor_cse_462 ^ state_4_3_31_0_sva_10 ^ state_2_10_1_lpi_4
      ^ plaintext_31_0_sva_10);
  assign xor_65_nl = state_2_4_1_lpi_6 ^ (key4[4]);
  assign state_xnor_165_nl = ~(xor_cse_465 ^ xor_cse_834 ^ xor_cse_842 ^ state_1_1_31_0_lpi_4_4
      ^ state_1_1_31_0_lpi_4_5);
  assign state_xnor_167_nl = ~(xor_cse_835 ^ xor_cse_1293 ^ plaintext_31_0_sva_5
      ^ plaintext_31_0_sva_6 ^ xor_cse_464 ^ state_4_3_31_0_sva_11 ^ state_2_11_1_lpi_4
      ^ plaintext_31_0_sva_11);
  assign xor_63_nl = state_2_5_1_lpi_6 ^ (key4[5]);
  assign state_xnor_168_nl = ~(xor_cse_466 ^ xor_cse_842 ^ state_1_1_31_0_lpi_4_5
      ^ Encrypt_Top_sbox_1_and_768 ^ state_4_4_6_lpi_3 ^ state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6])
      ^ state_1_1_31_0_lpi_4_6);
  assign state_xnor_170_nl = ~(xor_cse_1293 ^ xor_cse_1303 ^ plaintext_31_0_sva_6
      ^ plaintext_31_0_sva_7 ^ xor_cse_476 ^ state_4_3_31_0_sva_12 ^ state_2_12_1_lpi_4
      ^ plaintext_31_0_sva_12);
  assign xor_61_nl = state_2_6_1_lpi_6 ^ (key4[6]);
  assign state_xnor_171_nl = ~(xor_cse_477 ^ xor_cse_1306 ^ Encrypt_Top_sbox_1_and_768
      ^ state_4_4_6_lpi_3 ^ state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_71f1e461b47171ea32296c1ee9b3c00b2e_1[6])
      ^ state_1_1_31_0_lpi_4_6 ^ state_1_1_31_0_lpi_4_7);
  assign state_xnor_173_nl = ~(plaintext_31_0_sva_13 ^ xor_cse_1303 ^ xor_cse_845
      ^ plaintext_31_0_sva_7 ^ xor_cse_487 ^ state_4_3_31_0_sva_13 ^ state_2_13_1_lpi_4);
  assign xor_59_nl = state_2_7_1_lpi_6 ^ (key4[7]);
  assign state_xnor_174_nl = ~(state_1_1_63_32_lpi_4_8 ^ xor_cse_488 ^ xor_cse_1306
      ^ state_1_1_31_0_lpi_4_7 ^ Encrypt_Top_sbox_1_and_880 ^ state_4_4_8_lpi_3 ^
      state_2_8_1_lpi_4);
  assign ADLEN_i_ADLEN_i_mux_nl = MUX_v_4_2_2((z_out_2[3:0]), 4'b0001, fsm_output[8]);
  assign nor_28_nl = ~((ADLEN_i_7_0_sva_6_0_mx0c3 & (~ or_1265_cse)) | and_740_cse);
  assign state_xor_466_nl = xor_cse_2086 ^ Encrypt_Top_sbox_1_and_1_cse_0_sva_1 ^
      state_1_1_63_32_lpi_4_7 ^ xor_cse_196 ^ xor_cse_164 ^ xor_cse_2089 ^ xor_cse_2091
      ^ Encrypt_Top_sbox_1_and_628 ^ state_2_0_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]);
  assign state_xor_467_nl = xor_cse_2086 ^ Encrypt_Top_sbox_2_and_1_cse_0_sva_1 ^
      state_1_1_63_32_lpi_4_7 ^ xor_cse_196 ^ xor_cse_164 ^ xor_cse_2089 ^ xor_cse_2095
      ^ Encrypt_Top_sbox_1_and_628 ^ state_2_0_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]);
  assign xor_136_nl = state_1_1_31_0_lpi_4_0 ^ (key2[0]);
  assign state_xor_468_nl = xor_cse_2096 ^ xor_cse_2098 ^ xor_cse_2100 ^ Encrypt_Top_sbox_3_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1;
  assign state_xor_470_nl = xor_cse_2108 ^ xor_cse_2110 ^ xor_cse_2111;
  assign state_xor_471_nl = xor_cse_2114 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ Encrypt_Top_sbox_2_and_1_cse_1_sva_1 ^ xor_cse_2111;
  assign xor_134_nl = state_1_1_31_0_lpi_4_1 ^ (key2[1]);
  assign state_xor_472_nl = xor_cse_2118 ^ xor_cse_2120 ^ xor_cse_206 ^ xor_cse_2123
      ^ Encrypt_Top_sbox_1_and_630 ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1;
  assign state_xor_474_nl = xor_cse_2129 ^ xor_cse_185 ^ xor_cse_2131 ^ xor_cse_2132
      ^ xor_cse_2134 ^ state_2_2_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_2_sva_1;
  assign state_xor_475_nl = xor_cse_2129 ^ xor_cse_185 ^ xor_cse_2131 ^ xor_cse_2132
      ^ xor_cse_2137 ^ state_2_2_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_2_sva_1;
  assign xor_132_nl = state_1_1_31_0_lpi_4_2 ^ (key2[2]);
  assign state_xor_476_nl = xor_cse_2138 ^ Encrypt_Top_sbox_3_and_1_cse_41_sva_1
      ^ state_1_1_63_32_lpi_4_15 ^ xor_cse_217 ^ xor_cse_130 ^ xor_cse_2142 ^ Encrypt_Top_sbox_1_and_632
      ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1 ^ Encrypt_Top_sbox_1_and_588 ^ xor_cse_2145;
  assign state_xor_478_nl = xor_cse_2148 ^ xor_cse_2151 ^ xor_cse_2153 ^ state_2_3_1_lpi_4
      ^ Encrypt_Top_sbox_1_and_1_cse_3_sva_1 ^ xor_cse_2091 ^ state_2_0_1_lpi_4 ^
      Encrypt_Top_sbox_1_and_1_cse_0_sva_1;
  assign state_xor_479_nl = xor_cse_2148 ^ xor_cse_2151 ^ xor_cse_2157 ^ state_2_3_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_3_sva_1 ^ xor_cse_2095 ^ state_2_0_1_lpi_6 ^
      Encrypt_Top_sbox_2_and_1_cse_0_sva_1;
  assign xor_130_nl = state_1_1_31_0_lpi_4_3 ^ (key2[3]);
  assign state_xor_480_nl = xor_cse_2100 ^ xor_cse_2159 ^ xor_cse_228 ^ xor_cse_2162
      ^ Encrypt_Top_sbox_1_and_634 ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1;
  assign state_xor_482_nl = xor_cse_2167 ^ xor_cse_2168 ^ xor_cse_2109 ^ xor_cse_2172
      ^ state_2_4_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1 ^ xor_cse_2110;
  assign state_xor_483_nl = xor_cse_2167 ^ xor_cse_2168 ^ xor_cse_2115 ^ xor_cse_2176
      ^ state_2_4_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_4_sva_1 ^ state_2_1_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_1_sva_1;
  assign xor_128_nl = state_1_1_31_0_lpi_4_4 ^ (key2[4]);
  assign state_xor_484_nl = xor_cse_2178 ^ Encrypt_Top_sbox_1_and_636 ^ Encrypt_Top_sbox_1_and_630
      ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1 ^ xor_cse_238 ^ xor_cse_206 ^ xor_cse_2123
      ^ xor_cse_2182;
  assign state_xor_486_nl = xor_cse_2187 ^ state_2_2_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_2_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_44_sva_1 ^ xor_cse_217 ^ xor_cse_248 ^ xor_cse_2190
      ^ xor_cse_2192 ^ state_2_5_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_5_sva_1 ^
      xor_cse_2134;
  assign state_xor_487_nl = xor_cse_2187 ^ state_2_2_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_2_sva_1
      ^ Encrypt_Top_sbox_1_and_1_cse_44_sva_1 ^ xor_cse_217 ^ xor_cse_248 ^ xor_cse_2190
      ^ xor_cse_2196 ^ state_2_5_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_5_sva_1 ^
      xor_cse_2137;
  assign xor_126_nl = state_1_1_31_0_lpi_4_5 ^ (key2[5]);
  assign state_xor_488_nl = xor_cse_2197 ^ Encrypt_Top_sbox_1_and_632 ^ Encrypt_Top_sbox_1_and_576
      ^ xor_cse_2201 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1 ^ state_1_1_63_32_lpi_4_18
      ^ xor_cse_217 ^ xor_cse_35 ^ xor_cse_2142;
  assign state_xor_490_nl = xor_cse_2204 ^ xor_cse_2205 ^ xor_cse_2209 ^ state_2_6_1_lpi_4
      ^ Encrypt_Top_sbox_1_and_1_cse_6_sva_1 ^ xor_cse_2153 ^ state_2_3_1_lpi_4 ^
      Encrypt_Top_sbox_1_and_1_cse_3_sva_1;
  assign state_xor_491_nl = xor_cse_2204 ^ xor_cse_2205 ^ xor_cse_2213 ^ state_2_6_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_6_sva_1 ^ xor_cse_2157 ^ state_2_3_1_lpi_6 ^
      Encrypt_Top_sbox_2_and_1_cse_3_sva_1;
  assign xor_124_nl = state_1_1_31_0_lpi_4_6 ^ (key2[6]);
  assign state_xor_492_nl = xor_cse_2215 ^ Encrypt_Top_sbox_1_and_640 ^ Encrypt_Top_sbox_1_and_634
      ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1 ^ xor_cse_228 ^ xor_cse_258 ^ xor_cse_2162
      ^ xor_cse_2219;
  assign state_xor_494_nl = xor_cse_2224 ^ state_2_4_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1
      ^ state_1_1_63_32_lpi_4_14 ^ xor_cse_238 ^ xor_cse_268 ^ xor_cse_2227 ^ xor_cse_2229
      ^ state_2_7_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_7_sva_1 ^ xor_cse_2172;
  assign state_xor_495_nl = xor_cse_2224 ^ xor_cse_2230 ^ xor_cse_238 ^ xor_cse_2227
      ^ xor_cse_2176 ^ state_2_4_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_4_sva_1 ^
      state_1_1_63_32_lpi_4_14;
  assign xor_122_nl = state_1_1_31_0_lpi_4_7 ^ (key2[7]);
  assign state_xor_496_nl = xor_cse_2234 ^ xor_cse_2237 ^ xor_cse_238 ^ xor_cse_2182
      ^ Encrypt_Top_sbox_1_and_636 ^ Encrypt_Top_sbox_3_and_1_cse_46_sva_1;
  assign state_xor_498_nl = xor_cse_2242 ^ xor_cse_2243 ^ xor_cse_178 ^ xor_cse_2245
      ^ state_2_7_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_7_sva_1 ^ state_1_1_63_32_lpi_4_17;
  assign state_xor_499_nl = xor_cse_2242 ^ xor_cse_2230 ^ xor_cse_178 ^ xor_cse_2245
      ^ Encrypt_Top_sbox_1_and_642 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7])
      ^ state_1_1_63_32_lpi_4_17;
  assign xor_116_nl = state_1_1_31_0_lpi_4_10 ^ (key2[10]);
  assign state_xor_500_nl = xor_cse_2234 ^ xor_cse_2249 ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1
      ^ xor_cse_178 ^ xor_cse_2245;
  assign state_xor_544_nl = xor_cse_2388 ^ xor_cse_2389 ^ xor_cse_2091 ^ state_2_0_1_lpi_4
      ^ Encrypt_Top_sbox_1_and_1_cse_0_sva_1;
  assign state_xor_545_nl = xor_cse_2388 ^ xor_cse_2389 ^ xor_cse_2095 ^ state_2_0_1_lpi_6
      ^ Encrypt_Top_sbox_2_and_1_cse_0_sva_1;
  assign xor_86_nl = state_1_1_31_0_lpi_4_25 ^ (key2[25]);
  assign state_xor_546_nl = xor_cse_325 ^ xor_cse_2100 ^ xor_cse_2389;
  assign state_xor_548_nl = state_2_1_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_1_sva_1
      ^ xor_cse_2108 ^ xor_cse_2395;
  assign state_xor_549_nl = (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[1])
      ^ Encrypt_Top_sbox_2_and_1_cse_1_sva_1 ^ xor_cse_2395 ^ xor_cse_2114;
  assign xor_84_nl = state_1_1_31_0_lpi_4_26 ^ (key2[26]);
  assign state_xor_550_nl = Encrypt_Top_sbox_1_and_630 ^ xor_cse_206 ^ xor_cse_2123
      ^ xor_cse_2395;
  assign state_xor_552_nl = xor_cse_2399 ^ xor_cse_316 ^ xor_cse_2383 ^ xor_cse_2134
      ^ state_2_2_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2])
      ^ Encrypt_Top_sbox_1_and_1_cse_2_sva_1;
  assign state_xor_553_nl = xor_cse_2399 ^ xor_cse_316 ^ xor_cse_2383 ^ xor_cse_2137
      ^ state_2_2_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[2])
      ^ Encrypt_Top_sbox_2_and_1_cse_2_sva_1;
  assign xor_82_nl = state_1_1_31_0_lpi_4_27 ^ (key2[27]);
  assign state_xor_554_nl = xor_cse_316 ^ xor_cse_2142 ^ xor_cse_2383 ^ xor_cse_2399;
  assign state_xor_556_nl = xor_cse_2407 ^ xor_cse_325 ^ xor_cse_2390 ^ xor_cse_2153
      ^ state_2_3_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3])
      ^ Encrypt_Top_sbox_1_and_1_cse_3_sva_1;
  assign state_xor_557_nl = xor_cse_2407 ^ xor_cse_325 ^ xor_cse_2390 ^ xor_cse_2157
      ^ state_2_3_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[3])
      ^ Encrypt_Top_sbox_2_and_1_cse_3_sva_1;
  assign xor_80_nl = state_1_1_31_0_lpi_4_28 ^ (key2[28]);
  assign state_xor_558_nl = xor_cse_325 ^ xor_cse_2162 ^ xor_cse_2390 ^ xor_cse_2407;
  assign state_xor_560_nl = xor_cse_2414 ^ xor_cse_2396 ^ xor_cse_2416 ^ xor_cse_2172
      ^ state_2_4_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4])
      ^ Encrypt_Top_sbox_1_and_1_cse_4_sva_1;
  assign state_xor_561_nl = xor_cse_2414 ^ xor_cse_2396 ^ xor_cse_2416 ^ xor_cse_2176
      ^ state_2_4_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[4])
      ^ Encrypt_Top_sbox_2_and_1_cse_4_sva_1;
  assign xor_78_nl = state_1_1_31_0_lpi_4_29 ^ (key2[29]);
  assign state_xor_562_nl = xor_cse_2396 ^ xor_cse_2182 ^ xor_cse_2416 ^ xor_cse_2414;
  assign state_xor_564_nl = Encrypt_Top_sbox_1_and_638 ^ xor_cse_248 ^ xor_cse_343
      ^ xor_cse_384 ^ xor_cse_2400 ^ xor_cse_2422 ^ xor_cse_2423;
  assign state_xor_565_nl = Encrypt_Top_sbox_2_and_1_cse_5_sva_1 ^ xor_cse_248 ^
      xor_cse_343 ^ xor_cse_384 ^ xor_cse_2400 ^ xor_cse_2422 ^ xor_cse_2196 ^ Encrypt_Top_sbox_1_and_638
      ^ state_2_5_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5]);
  assign xor_76_nl = state_1_1_31_0_lpi_4_30 ^ (key2[30]);
  assign state_xor_566_nl = xor_cse_2197 ^ xor_cse_343 ^ xor_cse_384 ^ xor_cse_2400
      ^ xor_cse_2422;
  assign state_xor_568_nl = xor_cse_2427 ^ xor_cse_2408 ^ xor_cse_2429 ^ xor_cse_2209
      ^ state_2_6_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6])
      ^ Encrypt_Top_sbox_1_and_1_cse_6_sva_1;
  assign state_xor_569_nl = xor_cse_2427 ^ xor_cse_2408 ^ xor_cse_2429 ^ xor_cse_2213
      ^ state_2_6_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[6])
      ^ Encrypt_Top_sbox_2_and_1_cse_6_sva_1;
  assign xor_5_nl = state_1_1_31_0_lpi_4_31 ^ (key2[31]);
  assign state_xor_570_nl = xor_cse_2408 ^ xor_cse_2219 ^ xor_cse_2429 ^ xor_cse_2427;
  assign state_xor_502_nl = xor_cse_2255 ^ xor_cse_2256 ^ state_1_1_63_32_lpi_4_18
      ^ xor_cse_189 ^ xor_cse_278 ^ xor_cse_2258;
  assign xor_114_nl = state_1_1_31_0_lpi_4_11 ^ (key2[11]);
  assign state_xor_503_nl = xor_cse_2259 ^ xor_cse_2261 ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1
      ^ xor_cse_189 ^ xor_cse_278 ^ xor_cse_2258;
  assign state_xor_505_nl = xor_cse_2268 ^ xor_cse_2269 ^ state_1_1_63_32_lpi_4_19
      ^ xor_cse_204 ^ xor_cse_286 ^ xor_cse_2271;
  assign xor_112_nl = state_1_1_31_0_lpi_4_12 ^ (key2[12]);
  assign state_xor_506_nl = xor_cse_2272 ^ xor_cse_2274 ^ xor_cse_204 ^ xor_cse_2271
      ^ state_1_1_63_32_lpi_4_9 ^ Encrypt_Top_sbox_3_and_1_cse_51_sva_1;
  assign state_xor_508_nl = xor_cse_2280 ^ xor_cse_2281 ^ Encrypt_Top_sbox_1_and_1_cse_52_sva_1
      ^ xor_cse_178 ^ xor_cse_211 ^ xor_cse_2245;
  assign xor_110_nl = state_1_1_31_0_lpi_4_13 ^ (key2[13]);
  assign state_xor_509_nl = xor_cse_2280 ^ xor_cse_2283 ^ state_1_1_63_32_lpi_4_25
      ^ xor_cse_178 ^ xor_cse_211 ^ xor_cse_2245;
  assign state_xor_511_nl = xor_cse_2289 ^ xor_cse_2290 ^ xor_cse_189 ^ xor_cse_2258
      ^ Encrypt_Top_sbox_1_and_652 ^ Encrypt_Top_sbox_1_and_1_cse_53_sva_1;
  assign xor_108_nl = state_1_1_31_0_lpi_4_14 ^ (key2[14]);
  assign state_xor_512_nl = xor_cse_2289 ^ xor_cse_2293 ^ xor_cse_189 ^ xor_cse_2258
      ^ Encrypt_Top_sbox_1_and_652 ^ state_1_1_63_32_lpi_4_26;
  assign state_xor_514_nl = xor_cse_2298 ^ xor_cse_2299 ^ xor_cse_204 ^ xor_cse_2271
      ^ Encrypt_Top_sbox_1_and_654 ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1;
  assign xor_106_nl = state_1_1_31_0_lpi_4_15 ^ (key2[15]);
  assign state_xor_515_nl = xor_cse_2298 ^ xor_cse_2302 ^ xor_cse_204 ^ xor_cse_2271
      ^ Encrypt_Top_sbox_1_and_654 ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1;
  assign state_xor_517_nl = xor_cse_2308 ^ xor_cse_2309 ^ xor_cse_211 ^ xor_cse_2280
      ^ Encrypt_Top_sbox_1_and_656 ^ state_1_1_63_32_lpi_4_23;
  assign xor_104_nl = state_1_1_31_0_lpi_4_16 ^ (key2[16]);
  assign state_xor_518_nl = xor_cse_2308 ^ Encrypt_Top_sbox_1_and_656 ^ Encrypt_Top_sbox_1_and_532
      ^ xor_cse_2313 ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1 ^ state_1_1_63_32_lpi_4_28
      ^ xor_cse_211 ^ xor_cse_91 ^ xor_cse_2280;
  assign state_xor_520_nl = xor_cse_2289 ^ xor_cse_2319 ^ xor_cse_252 ^ xor_cse_2321
      ^ Encrypt_Top_sbox_1_and_652 ^ state_1_1_63_32_lpi_4_24;
  assign xor_102_nl = state_1_1_31_0_lpi_4_17 ^ (key2[17]);
  assign state_xor_521_nl = xor_cse_2289 ^ xor_cse_2323 ^ xor_cse_252 ^ xor_cse_2321
      ^ Encrypt_Top_sbox_1_and_652 ^ state_1_1_63_32_lpi_4_29;
  assign state_xor_523_nl = xor_cse_2298 ^ xor_cse_2330 ^ xor_cse_119 ^ xor_cse_2333;
  assign xor_100_nl = state_1_1_31_0_lpi_4_18 ^ (key2[18]);
  assign state_xor_524_nl = xor_cse_2298 ^ xor_cse_2330 ^ xor_cse_119 ^ xor_cse_2336
      ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1 ^ state_1_1_63_32_lpi_4_3;
  assign state_xor_526_nl = xor_cse_2308 ^ xor_cse_2340 ^ xor_cse_274 ^ xor_cse_2342
      ^ Encrypt_Top_sbox_1_and_656 ^ state_1_1_63_32_lpi_4_26;
  assign xor_98_nl = state_1_1_31_0_lpi_4_19 ^ (key2[19]);
  assign state_xor_527_nl = xor_cse_2308 ^ xor_cse_2344 ^ xor_cse_274 ^ xor_cse_2342
      ^ Encrypt_Top_sbox_1_and_656 ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1;
  assign state_xor_529_nl = xor_cse_2351 ^ xor_cse_2352 ^ xor_cse_252 ^ xor_cse_2321
      ^ Encrypt_Top_sbox_1_and_664 ^ state_1_1_63_32_lpi_4_27;
  assign xor_96_nl = state_1_1_31_0_lpi_4_20 ^ (key2[20]);
  assign state_xor_530_nl = xor_cse_2351 ^ Encrypt_Top_sbox_1_and_664 ^ Encrypt_Top_sbox_1_and_524
      ^ xor_cse_2356 ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1 ^ state_1_1_63_32_lpi_4_31
      ^ xor_cse_142 ^ xor_cse_252 ^ xor_cse_2321;
  assign state_xor_532_nl = xor_cse_2360 ^ xor_cse_2361 ^ xor_cse_2331 ^ Encrypt_Top_sbox_1_and_734
      ^ Encrypt_Top_sbox_1_and_1_cse_60_sva_1 ^ state_1_1_63_32_lpi_4_28;
  assign xor_94_nl = state_1_1_31_0_lpi_4_21 ^ (key2[21]);
  assign state_xor_533_nl = xor_cse_2360 ^ xor_cse_2361 ^ xor_cse_2331 ^ xor_cse_2366
      ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1 ^ state_1_1_63_32_lpi_4_4;
  assign state_xor_535_nl = xor_cse_164 ^ xor_cse_2089 ^ xor_cse_2371;
  assign xor_92_nl = state_1_1_31_0_lpi_4_22 ^ (key2[22]);
  assign state_xor_536_nl = Encrypt_Top_sbox_3_and_1_cse_61_sva_1 ^ xor_cse_2096
      ^ xor_cse_2371;
  assign state_xor_538_nl = xor_cse_2375 ^ xor_cse_2351 ^ Encrypt_Top_sbox_1_and_664
      ^ xor_cse_174 ^ xor_cse_308 ^ xor_cse_2112;
  assign xor_90_nl = state_1_1_31_0_lpi_4_23 ^ (key2[23]);
  assign state_xor_539_nl = xor_cse_2351 ^ xor_cse_2120 ^ xor_cse_308 ^ xor_cse_2375
      ^ Encrypt_Top_sbox_1_and_664 ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1;
  assign state_xor_541_nl = xor_cse_2132 ^ xor_cse_2360 ^ Encrypt_Top_sbox_1_and_666
      ^ xor_cse_185 ^ xor_cse_316 ^ xor_cse_2383;
  assign xor_88_nl = state_1_1_31_0_lpi_4_24 ^ (key2[24]);
  assign state_xor_542_nl = xor_cse_2360 ^ xor_cse_2138 ^ xor_cse_316 ^ xor_cse_2383
      ^ Encrypt_Top_sbox_1_and_666 ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1;
  assign state_xor_572_nl = xor_cse_2423 ^ xor_cse_2435 ^ xor_cse_2255 ^ xor_cse_2436;
  assign state_xor_573_nl = xor_cse_2436 ^ xor_cse_2435 ^ xor_cse_2255 ^ xor_cse_2196
      ^ state_2_5_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[5])
      ^ Encrypt_Top_sbox_2_and_1_cse_5_sva_1;
  assign xor_75_nl = state_1_1_63_32_lpi_4_0 ^ (key1[0]);
  assign state_xor_574_nl = xor_cse_2234 ^ xor_cse_2439 ^ Encrypt_Top_sbox_3_and_1_cse_32_sva_1
      ^ xor_cse_369 ^ xor_cse_2416;
  assign state_xor_575_nl = xor_cse_2442 ^ xor_cse_2443 ^ xor_cse_286 ^ xor_cse_2268
      ^ xor_cse_2209 ^ state_2_6_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_6_sva_1;
  assign state_xor_576_nl = xor_cse_2442 ^ xor_cse_2443 ^ xor_cse_286 ^ xor_cse_2268
      ^ xor_cse_2213 ^ state_2_6_1_lpi_6 ^ Encrypt_Top_sbox_2_and_1_cse_6_sva_1;
  assign xor_77_nl = state_1_1_63_32_lpi_4_1 ^ (key1[1]);
  assign state_xor_577_nl = xor_cse_2448 ^ Encrypt_Top_sbox_1_and_620 ^ Encrypt_Top_sbox_1_and_534
      ^ xor_cse_2262 ^ Encrypt_Top_sbox_3_and_1_cse_8_sva_1 ^ state_1_1_63_32_lpi_4_8
      ^ xor_cse_278 ^ xor_cse_384 ^ xor_cse_2422;
  assign state_xor_578_nl = xor_cse_2452 ^ xor_cse_2243 ^ xor_cse_369 ^ xor_cse_2416
      ^ state_1_1_63_32_lpi_4_0 ^ state_2_7_1_lpi_4 ^ Encrypt_Top_sbox_1_and_1_cse_7_sva_1;
  assign state_xor_579_nl = xor_cse_2452 ^ xor_cse_2230 ^ xor_cse_369 ^ xor_cse_2416
      ^ state_1_1_63_32_lpi_4_0 ^ Encrypt_Top_sbox_1_and_642 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]);
  assign xor_79_nl = state_1_1_63_32_lpi_4_2 ^ (key1[2]);
  assign state_xor_580_nl = xor_cse_2457 ^ xor_cse_2274 ^ xor_cse_394 ^ xor_cse_2429
      ^ state_1_1_63_32_lpi_4_0 ^ state_1_1_63_32_lpi_4_9;
  assign state_xor_581_nl = xor_cse_2255 ^ xor_cse_2461 ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1
      ^ xor_cse_278 ^ xor_cse_384 ^ xor_cse_2422;
  assign xor_81_nl = state_1_1_63_32_lpi_4_3 ^ (key1[3]);
  assign state_xor_582_nl = xor_cse_2463 ^ xor_cse_2439 ^ xor_cse_178 ^ xor_cse_2245
      ^ state_1_1_63_32_lpi_4_1 ^ Encrypt_Top_sbox_3_and_1_cse_32_sva_1;
  assign state_xor_583_nl = xor_cse_2151 ^ xor_cse_2086 ^ state_1_1_63_32_lpi_4_7
      ^ xor_cse_252 ^ xor_cse_8 ^ xor_cse_2321;
  assign xor_83_nl = state_1_1_63_32_lpi_4_4 ^ (key1[4]);
  assign state_xor_584_nl = xor_cse_2468 ^ xor_cse_2448 ^ xor_cse_2469;
  assign state_xor_585_nl = xor_cse_2331 ^ xor_cse_2167 ^ state_1_1_63_32_lpi_4_11
      ^ xor_cse_263 ^ xor_cse_120 ^ xor_cse_2113;
  assign xor_85_nl = state_1_1_63_32_lpi_4_5 ^ (key1[5]);
  assign state_xor_586_nl = xor_cse_2472 ^ xor_cse_2457 ^ xor_cse_204 ^ xor_cse_2271
      ^ state_1_1_63_32_lpi_4_11 ^ state_1_1_63_32_lpi_4_0;
  assign state_xor_587_nl = Encrypt_Top_sbox_1_and_1_cse_44_sva_1 ^ xor_cse_2131
      ^ xor_cse_2187 ^ xor_cse_2476;
  assign xor_87_nl = state_1_1_63_32_lpi_4_6 ^ (key1[6]);
  assign state_xor_588_nl = xor_cse_2463 ^ xor_cse_2477 ^ xor_cse_211 ^ xor_cse_2280
      ^ state_1_1_63_32_lpi_4_12 ^ state_1_1_63_32_lpi_4_1;
  assign state_xor_589_nl = xor_cse_2351 ^ xor_cse_2204 ^ xor_cse_8 ^ xor_cse_2151
      ^ state_1_1_63_32_lpi_4_13 ^ Encrypt_Top_sbox_1_and_664;
  assign xor_89_nl = state_1_1_63_32_lpi_4_7 ^ (key1[7]);
  assign state_xor_590_nl = xor_cse_2289 ^ xor_cse_2469 ^ xor_cse_2098 ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1
      ^ Encrypt_Top_sbox_1_and_608 ^ Encrypt_Top_sbox_1_and_652;
  assign state_xor_591_nl = xor_cse_2360 ^ xor_cse_2167 ^ xor_cse_2224 ^ state_1_1_63_32_lpi_4_14
      ^ state_1_1_63_32_lpi_4_11 ^ Encrypt_Top_sbox_1_and_666;
  assign xor_91_nl = state_1_1_63_32_lpi_4_8 ^ (key1[8]);
  assign state_xor_592_nl = xor_cse_2298 ^ xor_cse_2472 ^ xor_cse_2118 ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1
      ^ state_1_1_63_32_lpi_4_11 ^ Encrypt_Top_sbox_1_and_654;
  assign state_xor_593_nl = xor_cse_2435 ^ xor_cse_2187 ^ Encrypt_Top_sbox_1_and_1_cse_44_sva_1
      ^ xor_cse_77 ^ xor_cse_299 ^ xor_cse_2372;
  assign xor_93_nl = state_1_1_63_32_lpi_4_9 ^ (key1[9]);
  assign state_xor_594_nl = xor_cse_2308 ^ xor_cse_2477 ^ xor_cse_130 ^ xor_cse_2488
      ^ state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_1_and_656;
  assign state_xor_595_nl = xor_cse_2204 ^ xor_cse_2443 ^ xor_cse_308 ^ xor_cse_2375
      ^ Encrypt_Top_sbox_1_and_560 ^ state_1_1_63_32_lpi_4_13;
  assign xor_95_nl = state_1_1_63_32_lpi_4_10 ^ (key1[10]);
  assign state_xor_596_nl = xor_cse_2098 ^ xor_cse_2159 ^ xor_cse_252 ^ xor_cse_2321
      ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_39_sva_1;
  assign state_xor_597_nl = xor_cse_2242 ^ xor_cse_2224 ^ xor_cse_316 ^ xor_cse_2383
      ^ state_1_1_63_32_lpi_4_17 ^ state_1_1_63_32_lpi_4_14;
  assign xor_97_nl = state_1_1_63_32_lpi_4_11 ^ (key1[11]);
  assign state_xor_598_nl = xor_cse_2118 ^ xor_cse_2178 ^ xor_cse_263 ^ xor_cse_2331
      ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_40_sva_1;
  assign state_xor_599_nl = xor_cse_2435 ^ xor_cse_2256 ^ state_1_1_63_32_lpi_4_18
      ^ xor_cse_77 ^ xor_cse_325 ^ xor_cse_2390;
  assign xor_99_nl = state_1_1_63_32_lpi_4_12 ^ (key1[12]);
  assign state_xor_600_nl = xor_cse_2476 ^ xor_cse_35 ^ Encrypt_Top_sbox_1_and_576
      ^ xor_cse_2201 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1 ^ state_1_1_63_32_lpi_4_18
      ^ xor_cse_2488;
  assign state_xor_601_nl = xor_cse_2269 ^ xor_cse_2443 ^ xor_cse_334 ^ xor_cse_2396
      ^ state_1_1_63_32_lpi_4_19 ^ Encrypt_Top_sbox_1_and_560;
  assign xor_101_nl = state_1_1_63_32_lpi_4_13 ^ (key1[13]);
  assign state_xor_602_nl = xor_cse_2351 ^ xor_cse_2215 ^ xor_cse_2159 ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_42_sva_1 ^ Encrypt_Top_sbox_1_and_664;
  assign state_xor_603_nl = xor_cse_2268 ^ xor_cse_2505 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1
      ^ xor_cse_286 ^ xor_cse_394 ^ xor_cse_2429;
  assign xor_103_nl = state_1_1_63_32_lpi_4_14 ^ (key1[14]);
  assign state_xor_604_nl = xor_cse_2360 ^ xor_cse_2237 ^ xor_cse_2178 ^ Encrypt_Top_sbox_3_and_1_cse_46_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_43_sva_1 ^ Encrypt_Top_sbox_1_and_666;
  assign state_xor_605_nl = xor_cse_2242 ^ xor_cse_2281 ^ xor_cse_343 ^ xor_cse_2400
      ^ Encrypt_Top_sbox_1_and_1_cse_52_sva_1 ^ state_1_1_63_32_lpi_4_17;
  assign xor_105_nl = state_1_1_63_32_lpi_4_15 ^ (key1[15]);
  assign state_xor_606_nl = xor_cse_2510 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1
      ^ Encrypt_Top_sbox_1_and_576 ^ xor_cse_2201 ^ Encrypt_Top_sbox_3_and_1_cse_44_sva_1
      ^ state_1_1_63_32_lpi_4_18 ^ xor_cse_35 ^ xor_cse_299 ^ xor_cse_2372;
  assign state_xor_607_nl = xor_cse_2256 ^ xor_cse_2290 ^ xor_cse_357 ^ xor_cse_2408
      ^ Encrypt_Top_sbox_1_and_1_cse_53_sva_1 ^ state_1_1_63_32_lpi_4_18;
  assign xor_107_nl = state_1_1_63_32_lpi_4_16 ^ (key1[16]);
  assign state_xor_608_nl = xor_cse_2516 ^ xor_cse_2215 ^ xor_cse_308 ^ xor_cse_2375
      ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_45_sva_1;
  assign state_xor_609_nl = xor_cse_2269 ^ xor_cse_2299 ^ xor_cse_369 ^ xor_cse_2416
      ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1 ^ state_1_1_63_32_lpi_4_19;
  assign xor_109_nl = state_1_1_63_32_lpi_4_17 ^ (key1[17]);
  assign state_xor_610_nl = xor_cse_2237 ^ xor_cse_2249 ^ xor_cse_316 ^ xor_cse_2383
      ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_46_sva_1;
  assign state_xor_611_nl = xor_cse_2309 ^ xor_cse_2281 ^ xor_cse_384 ^ xor_cse_2422
      ^ state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_1_and_1_cse_52_sva_1;
  assign xor_111_nl = state_1_1_63_32_lpi_4_18 ^ (key1[18]);
  assign state_xor_612_nl = xor_cse_2510 ^ xor_cse_2259 ^ xor_cse_325 ^ xor_cse_2390
      ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1;
  assign state_xor_613_nl = xor_cse_2319 ^ xor_cse_2290 ^ xor_cse_394 ^ xor_cse_2429
      ^ state_1_1_63_32_lpi_4_24 ^ Encrypt_Top_sbox_1_and_1_cse_53_sva_1;
  assign xor_113_nl = state_1_1_63_32_lpi_4_19 ^ (key1[19]);
  assign state_xor_614_nl = xor_cse_2272 ^ xor_cse_2516 ^ xor_cse_334 ^ xor_cse_2396
      ^ Encrypt_Top_sbox_3_and_1_cse_51_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1;
  assign state_xor_615_nl = xor_cse_2452 ^ xor_cse_2299 ^ xor_cse_119 ^ Encrypt_Top_sbox_1_and_528
      ^ Encrypt_Top_sbox_1_and_728 ^ Encrypt_Top_sbox_1_and_1_cse_57_sva_1 ^ state_1_1_63_32_lpi_4_25
      ^ Encrypt_Top_sbox_1_and_1_cse_54_sva_1 ^ state_1_1_63_32_lpi_4_0;
  assign xor_115_nl = state_1_1_63_32_lpi_4_20 ^ (key1[20]);
  assign state_xor_616_nl = xor_cse_2283 ^ xor_cse_2249 ^ xor_cse_343 ^ xor_cse_2400
      ^ state_1_1_63_32_lpi_4_25 ^ Encrypt_Top_sbox_3_and_1_cse_49_sva_1;
  assign state_xor_617_nl = xor_cse_2309 ^ xor_cse_2340 ^ xor_cse_2461 ^ state_1_1_63_32_lpi_4_26
      ^ state_1_1_63_32_lpi_4_23 ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1;
  assign xor_117_nl = state_1_1_63_32_lpi_4_21 ^ (key1[21]);
  assign state_xor_618_nl = xor_cse_2293 ^ xor_cse_2259 ^ xor_cse_357 ^ xor_cse_2408
      ^ state_1_1_63_32_lpi_4_26 ^ Encrypt_Top_sbox_3_and_1_cse_50_sva_1;
  assign state_xor_619_nl = xor_cse_2352 ^ xor_cse_2319 ^ xor_cse_2505 ^ state_1_1_63_32_lpi_4_27
      ^ state_1_1_63_32_lpi_4_24 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1;
  assign xor_119_nl = state_1_1_63_32_lpi_4_22 ^ (key1[22]);
  assign state_xor_620_nl = xor_cse_2272 ^ xor_cse_2302 ^ xor_cse_369 ^ xor_cse_2416
      ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_51_sva_1;
  assign state_xor_621_nl = xor_cse_2543 ^ xor_cse_2544 ^ xor_cse_2545 ^ xor_cse_2333;
  assign xor_121_nl = state_1_1_63_32_lpi_4_23 ^ (key1[23]);
  assign state_xor_622_nl = xor_cse_2283 ^ Encrypt_Top_sbox_1_and_532 ^ xor_cse_2313
      ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1 ^ state_1_1_63_32_lpi_4_28 ^ state_1_1_63_32_lpi_4_25
      ^ xor_cse_91 ^ xor_cse_384 ^ xor_cse_2422;
  assign state_xor_623_nl = xor_cse_2340 ^ xor_cse_2549 ^ xor_cse_164 ^ xor_cse_2089
      ^ state_1_1_63_32_lpi_4_26 ^ Encrypt_Top_sbox_1_and_608;
  assign xor_123_nl = state_1_1_63_32_lpi_4_24 ^ (key1[24]);
  assign state_xor_624_nl = xor_cse_2293 ^ xor_cse_2323 ^ xor_cse_394 ^ xor_cse_2429
      ^ state_1_1_63_32_lpi_4_29 ^ state_1_1_63_32_lpi_4_26;
  assign state_xor_625_nl = xor_cse_2452 ^ xor_cse_2544 ^ xor_cse_178 ^ xor_cse_2245
      ^ state_1_1_63_32_lpi_4_3 ^ state_1_1_63_32_lpi_4_0;
  assign xor_125_nl = state_1_1_63_32_lpi_4_25 ^ (key1[25]);
  assign state_xor_626_nl = xor_cse_2302 ^ xor_cse_2439 ^ xor_cse_119 ^ Encrypt_Top_sbox_1_and_528
      ^ xor_cse_2336 ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1 ^ state_1_1_63_32_lpi_4_3
      ^ Encrypt_Top_sbox_3_and_1_cse_54_sva_1 ^ Encrypt_Top_sbox_3_and_1_cse_32_sva_1;
  assign state_xor_627_nl = xor_cse_2352 ^ xor_cse_2559 ^ xor_cse_174 ^ xor_cse_2112
      ^ state_1_1_63_32_lpi_4_27 ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1;
  assign xor_127_nl = state_1_1_63_32_lpi_4_26 ^ (key1[26]);
  assign state_xor_628_nl = xor_cse_2344 ^ xor_cse_2448 ^ xor_cse_91 ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1
      ^ Encrypt_Top_sbox_1_and_532 ^ xor_cse_2313 ^ Encrypt_Top_sbox_3_and_1_cse_55_sva_1
      ^ state_1_1_63_32_lpi_4_28 ^ Encrypt_Top_sbox_1_and_620;
  assign state_xor_629_nl = xor_cse_2565 ^ xor_cse_2545 ^ xor_cse_185 ^ xor_cse_2132
      ^ Encrypt_Top_sbox_1_and_522 ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1;
  assign xor_129_nl = state_1_1_63_32_lpi_4_27 ^ (key1[27]);
  assign state_xor_630_nl = xor_cse_2457 ^ xor_cse_2323 ^ xor_cse_142 ^ Encrypt_Top_sbox_1_and_524
      ^ xor_cse_2356 ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1 ^ state_1_1_63_32_lpi_4_31
      ^ state_1_1_63_32_lpi_4_29 ^ state_1_1_63_32_lpi_4_0;
  assign state_xor_631_nl = xor_cse_2468 ^ xor_cse_2549 ^ xor_cse_25 ^ Encrypt_Top_sbox_1_and_694
      ^ Encrypt_Top_sbox_1_and_1_cse_33_sva_1 ^ state_1_1_63_32_lpi_4_1;
  assign xor_131_nl = state_1_1_63_32_lpi_4_28 ^ (key1[28]);
  assign state_xor_632_nl = xor_cse_2543 ^ xor_cse_2463 ^ xor_cse_154 ^ xor_cse_2366
      ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1 ^ state_1_1_63_32_lpi_4_4 ^ xor_cse_2336
      ^ Encrypt_Top_sbox_3_and_1_cse_57_sva_1 ^ state_1_1_63_32_lpi_4_1;
  assign state_xor_633_nl = xor_cse_2505 ^ xor_cse_2559 ^ xor_cse_204 ^ xor_cse_2271
      ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_1_and_1_cse_34_sva_1;
  assign xor_133_nl = state_1_1_63_32_lpi_4_29 ^ (key1[29]);
  assign state_xor_634_nl = xor_cse_2096 ^ xor_cse_2344 ^ xor_cse_2469 ^ Encrypt_Top_sbox_3_and_1_cse_61_sva_1
      ^ Encrypt_Top_sbox_3_and_1_cse_58_sva_1 ^ Encrypt_Top_sbox_1_and_608;
  assign state_xor_635_nl = xor_cse_2565 ^ xor_cse_2544 ^ xor_cse_211 ^ xor_cse_2280
      ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1 ^ state_1_1_63_32_lpi_4_3;
  assign xor_135_nl = state_1_1_63_32_lpi_4_30 ^ (key1[30]);
  assign state_xor_636_nl = xor_cse_2472 ^ xor_cse_2120 ^ xor_cse_142 ^ Encrypt_Top_sbox_3_and_1_cse_62_sva_1
      ^ Encrypt_Top_sbox_1_and_524 ^ xor_cse_2356 ^ Encrypt_Top_sbox_3_and_1_cse_59_sva_1
      ^ state_1_1_63_32_lpi_4_31 ^ state_1_1_63_32_lpi_4_11;
  assign state_xor_637_nl = xor_cse_2289 ^ xor_cse_2086 ^ xor_cse_2549 ^ state_1_1_63_32_lpi_4_7
      ^ Encrypt_Top_sbox_1_and_608 ^ Encrypt_Top_sbox_1_and_652;
  assign xor_137_nl = state_1_1_63_32_lpi_4_31 ^ (key1[31]);
  assign state_xor_638_nl = xor_cse_2138 ^ xor_cse_2477 ^ xor_cse_154 ^ Encrypt_Top_sbox_3_and_1_cse_63_sva_1
      ^ Encrypt_Top_sbox_1_and_522 ^ xor_cse_2366 ^ Encrypt_Top_sbox_3_and_1_cse_60_sva_1
      ^ state_1_1_63_32_lpi_4_4 ^ state_1_1_63_32_lpi_4_12;
  assign state_xor_639_nl = xor_cse_2298 ^ xor_cse_2559 ^ xor_cse_120 ^ xor_cse_2113
      ^ Encrypt_Top_sbox_1_and_1_cse_37_sva_1 ^ Encrypt_Top_sbox_1_and_654;
  assign xor_120_nl = state_1_1_31_0_lpi_4_8 ^ (key2[8]);
  assign state_xor_640_nl = xor_cse_2510 ^ xor_cse_2197 ^ Encrypt_Top_sbox_3_and_1_cse_47_sva_1
      ^ xor_cse_278 ^ xor_cse_2261;
  assign state_xor_641_nl = xor_cse_2308 ^ xor_cse_2565 ^ xor_cse_130 ^ xor_cse_2131
      ^ Encrypt_Top_sbox_1_and_1_cse_38_sva_1 ^ Encrypt_Top_sbox_1_and_656;
  assign xor_118_nl = state_1_1_31_0_lpi_4_9 ^ (key2[9]);
  assign state_xor_642_nl = xor_cse_2516 ^ xor_cse_2274 ^ xor_cse_258 ^ xor_cse_2219
      ^ state_1_1_63_32_lpi_4_9 ^ Encrypt_Top_sbox_1_and_640 ^ Encrypt_Top_sbox_3_and_1_cse_48_sva_1;
  assign state_xor_643_nl = xor_cse_1845 ^ xor_cse_352 ^ xor_cse_933 ^ xor_cse_1849
      ^ (key2[0]) ^ xor_cse_1853 ^ xor_cse_1854 ^ state_4_3_31_0_sva_17;
  assign state_xor_644_nl = xor_cse_252 ^ xor_cse_1299 ^ xor_cse_2598 ^ xor_cse_1300;
  assign state_xor_645_nl = xor_cse_1300 ^ xor_cse_252 ^ xor_cse_1299 ^ Encrypt_Top_sbox_2_and_520
      ^ Encrypt_Top_sbox_2_and_522 ^ state_2_0_1_lpi_6 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[0]);
  assign state_xor_646_nl = xor_cse_1868 ^ xor_cse_1871 ^ (key2[1]) ^ xor_cse_364
      ^ xor_cse_1865;
  assign state_xor_647_nl = xor_cse_206 ^ xor_cse_189 ^ xor_cse_263 ^ xor_cse_1309
      ^ xor_cse_2602 ^ xor_cse_1310;
  assign state_xor_648_nl = xor_cse_2604 ^ xor_cse_189 ^ xor_cse_263 ^ xor_cse_1309
      ^ Encrypt_Top_sbox_2_and_530 ^ Encrypt_Top_sbox_2_and_610 ^ state_4_4_11_lpi_3;
  assign state_xor_649_nl = xor_cse_1886 ^ xor_cse_1889 ^ (key2[2]) ^ xor_cse_377
      ^ xor_cse_1883;
  assign state_xor_650_nl = state_2_2_1_lpi_4 ^ xor_cse_2278 ^ xor_cse_2608 ^ xor_cse_2279;
  assign state_xor_651_nl = state_2_2_1_lpi_6 ^ xor_cse_2278 ^ xor_cse_2608 ^ xor_cse_2279;
  assign state_xor_652_nl = xor_cse_1895 ^ xor_cse_1904 ^ (key2[3]) ^ xor_cse_389
      ^ xor_cse_1901;
  assign state_xor_653_nl = state_2_3_1_lpi_4 ^ xor_cse_2373 ^ xor_cse_2610 ^ xor_cse_2374;
  assign state_xor_654_nl = state_2_3_1_lpi_6 ^ xor_cse_2373 ^ xor_cse_2610 ^ xor_cse_2374;
  assign state_xor_655_nl = xor_cse_1877 ^ xor_cse_1916 ^ (key2[4]) ^ xor_cse_405
      ^ xor_cse_1913;
  assign state_xor_656_nl = xor_cse_2612 ^ xor_cse_221 ^ xor_cse_290 ^ xor_cse_2393
      ^ state_2_4_1_lpi_4 ^ Encrypt_Top_sbox_2_and_634 ^ state_4_4_14_lpi_3;
  assign state_xor_657_nl = xor_cse_2612 ^ xor_cse_221 ^ xor_cse_290 ^ xor_cse_2393
      ^ state_2_4_1_lpi_6 ^ Encrypt_Top_sbox_2_and_634 ^ state_4_4_14_lpi_3;
  assign state_xor_658_nl = xor_cse_1855 ^ xor_cse_1922 ^ (key2[5]) ^ xor_cse_417
      ^ xor_cse_1907;
  assign state_xor_659_nl = state_2_5_1_lpi_4 ^ xor_cse_2397 ^ xor_cse_2618 ^ xor_cse_2398;
  assign state_xor_660_nl = state_2_5_1_lpi_6 ^ xor_cse_2397 ^ xor_cse_2618 ^ xor_cse_2398;
  assign state_xor_661_nl = xor_cse_1835 ^ xor_cse_1928 ^ (key2[6]) ^ xor_cse_430
      ^ xor_cse_1892;
  assign state_xor_662_nl = state_2_6_1_lpi_4 ^ xor_cse_2405 ^ xor_cse_2620 ^ xor_cse_2406;
  assign state_xor_663_nl = state_2_6_1_lpi_6 ^ xor_cse_2405 ^ xor_cse_2620 ^ xor_cse_2406;
  assign state_xor_664_nl = xor_cse_1936 ^ xor_cse_444 ^ xor_cse_933 ^ xor_cse_1874
      ^ (key2[7]) ^ xor_cse_1853 ^ xor_cse_1854 ^ state_4_3_31_0_sva_17;
  assign state_xor_665_nl = xor_cse_1350 ^ xor_cse_2413 ^ xor_cse_268 ^ Encrypt_Top_sbox_2_and_576
      ^ Encrypt_Top_sbox_2_and_578 ^ state_2_7_1_lpi_4 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7]);
  assign state_xor_666_nl = xor_cse_268 ^ xor_cse_2625 ^ xor_cse_1350 ^ xor_cse_2413;
  assign state_xor_769_nl = xor_cse_1925 ^ xor_cse_1998 ^ (key1[15]) ^ xor_cse_352
      ^ xor_cse_1849;
  assign state_xor_770_nl = xor_cse_194 ^ xor_cse_196 ^ xor_cse_77 ^ xor_cse_2598
      ^ Encrypt_Top_sbox_2_and_646 ^ state_1_1_63_32_lpi_4_15 ^ state_1_1_63_32_lpi_4_25;
  assign state_xor_771_nl = xor_cse_194 ^ xor_cse_2808 ^ xor_cse_77 ^ Encrypt_Top_sbox_2_and_646
      ^ state_1_1_63_32_lpi_4_15 ^ state_1_1_63_32_lpi_4_25 ^ Encrypt_Top_sbox_2_and_522;
  assign state_xor_772_nl = state_1_1_63_32_lpi_4_3 ^ xor_cse_77 ^ xor_cse_194 ^
      xor_cse_195;
  assign state_xor_773_nl = xor_cse_1919 ^ xor_cse_1991 ^ (key1[16]) ^ xor_cse_364
      ^ xor_cse_1865;
  assign state_xor_774_nl = xor_cse_206 ^ xor_cse_2602 ^ xor_cse_2707 ^ xor_cse_2771;
  assign state_xor_775_nl = Encrypt_Top_sbox_2_and_530 ^ xor_cse_2707 ^ xor_cse_2771
      ^ xor_cse_2604;
  assign state_xor_776_nl = xor_cse_132 ^ xor_cse_94 ^ xor_cse_209 ^ xor_cse_205;
  assign state_xor_777_nl = xor_cse_1910 ^ xor_cse_1985 ^ (key1[17]) ^ xor_cse_377
      ^ xor_cse_1883;
  assign state_xor_778_nl = xor_cse_2608 ^ xor_cse_142 ^ xor_cse_10 ^ xor_cse_2814
      ^ Encrypt_Top_sbox_2_and_550 ^ state_1_1_63_32_lpi_4_27 ^ state_2_2_1_lpi_4;
  assign state_xor_779_nl = xor_cse_2608 ^ xor_cse_142 ^ xor_cse_10 ^ xor_cse_2814
      ^ Encrypt_Top_sbox_2_and_550 ^ state_1_1_63_32_lpi_4_27 ^ state_2_2_1_lpi_6;
  assign state_xor_780_nl = xor_cse_141 ^ xor_cse_217 ^ xor_cse_10 ^ xor_cse_218
      ^ Encrypt_Top_sbox_2_and_628 ^ Encrypt_Top_sbox_2_and_630 ^ state_1_1_63_32_lpi_4_22;
  assign state_xor_781_nl = xor_cse_1979 ^ xor_cse_1898 ^ (key1[18]) ^ xor_cse_389
      ^ xor_cse_1901;
  assign state_xor_782_nl = xor_cse_2610 ^ xor_cse_154 ^ xor_cse_24 ^ xor_cse_2822
      ^ Encrypt_Top_sbox_2_and_622 ^ state_1_1_63_32_lpi_4_18 ^ state_2_3_1_lpi_4;
  assign state_xor_783_nl = xor_cse_2610 ^ xor_cse_154 ^ xor_cse_24 ^ xor_cse_2822
      ^ Encrypt_Top_sbox_2_and_622 ^ state_1_1_63_32_lpi_4_18 ^ state_2_3_1_lpi_6;
  assign state_xor_784_nl = xor_cse_228 ^ xor_cse_229 ^ xor_cse_153 ^ xor_cse_226;
  assign state_xor_785_nl = xor_cse_1973 ^ xor_cse_1880 ^ (key1[19]) ^ xor_cse_405
      ^ xor_cse_1913;
  assign state_xor_786_nl = state_2_4_1_lpi_4 ^ xor_cse_236 ^ xor_cse_2612 ^ xor_cse_2827;
  assign state_xor_787_nl = state_2_4_1_lpi_6 ^ xor_cse_236 ^ xor_cse_2612 ^ xor_cse_2827;
  assign state_xor_788_nl = state_1_1_63_32_lpi_4_5 ^ xor_cse_238 ^ xor_cse_239 ^
      xor_cse_235;
  assign state_xor_789_nl = xor_cse_1966 ^ xor_cse_1969 ^ (key1[20]) ^ xor_cse_417
      ^ xor_cse_1907;
  assign state_xor_790_nl = xor_cse_2618 ^ xor_cse_2791 ^ state_2_5_1_lpi_4 ^ xor_cse_51
      ^ xor_cse_2830;
  assign state_xor_791_nl = xor_cse_2618 ^ xor_cse_2791 ^ state_2_5_1_lpi_6 ^ xor_cse_51
      ^ xor_cse_2830;
  assign state_xor_792_nl = xor_cse_246 ^ xor_cse_248 ^ xor_cse_51 ^ xor_cse_249
      ^ Encrypt_Top_sbox_2_and_606 ^ state_1_1_63_32_lpi_4_25 ^ state_1_1_63_32_lpi_4_6;
  assign state_xor_793_nl = xor_cse_1838 ^ xor_cse_1960 ^ (key1[21]) ^ xor_cse_430
      ^ xor_cse_1892;
  assign state_xor_794_nl = xor_cse_256 ^ xor_cse_258 ^ xor_cse_185 ^ xor_cse_2836
      ^ state_1_1_63_32_lpi_4_21 ^ state_1_1_63_32_lpi_4_31 ^ state_2_6_1_lpi_4;
  assign state_xor_795_nl = xor_cse_256 ^ xor_cse_258 ^ xor_cse_185 ^ xor_cse_2836
      ^ state_1_1_63_32_lpi_4_21 ^ state_1_1_63_32_lpi_4_31 ^ state_2_6_1_lpi_6;
  assign state_xor_796_nl = state_1_1_63_32_lpi_4_7 ^ xor_cse_260 ^ xor_cse_256 ^
      xor_cse_257;
  assign state_xor_797_nl = xor_cse_1874 ^ xor_cse_1951 ^ (key1[22]) ^ xor_cse_352
      ^ xor_cse_444 ^ xor_cse_1849;
  assign state_xor_798_nl = xor_cse_267 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7])
      ^ xor_cse_196 ^ xor_cse_2598 ^ state_1_1_63_32_lpi_4_22 ^ Encrypt_Top_sbox_2_and_576
      ^ Encrypt_Top_sbox_2_and_578 ^ state_2_7_1_lpi_4;
  assign state_xor_799_nl = xor_cse_267 ^ xor_cse_2808 ^ xor_cse_2625 ^ state_1_1_63_32_lpi_4_22
      ^ Encrypt_Top_sbox_2_and_522;
  assign state_xor_800_nl = xor_cse_267 ^ state_1_1_63_32_lpi_4_27 ^ xor_cse_196
      ^ xor_cse_197 ^ xor_cse_270;
  assign state_xor_801_nl = xor_cse_1941 ^ xor_cse_364 ^ xor_cse_1162 ^ xor_cse_1865
      ^ xor_cse_1862 ^ xor_cse_1864 ^ state_4_3_31_0_sva_8 ^ (key1[23]);
  assign state_xor_802_nl = xor_cse_206 ^ xor_cse_91 ^ xor_cse_278 ^ xor_cse_2602
      ^ xor_cse_2848 ^ Encrypt_Top_sbox_2_and_586 ^ state_1_1_31_0_lpi_4_8;
  assign state_xor_803_nl = xor_cse_2604 ^ xor_cse_91 ^ xor_cse_278 ^ xor_cse_2848
      ^ Encrypt_Top_sbox_2_and_530 ^ Encrypt_Top_sbox_2_and_586 ^ state_1_1_31_0_lpi_4_8;
  assign state_xor_804_nl = xor_cse_206 ^ xor_cse_207 ^ xor_cse_277 ^ xor_cse_172;
  assign state_xor_805_nl = xor_cse_1931 ^ xor_cse_377 ^ xor_cse_1172 ^ xor_cse_1883
      ^ xor_cse_1843 ^ xor_cse_1844 ^ state_4_3_31_0_sva_9 ^ (key1[24]);
  assign state_xor_806_nl = xor_cse_2608 ^ xor_cse_106 ^ xor_cse_286 ^ xor_cse_2855
      ^ Encrypt_Top_sbox_2_and_574 ^ state_1_1_63_32_lpi_4_24 ^ state_2_2_1_lpi_4;
  assign state_xor_807_nl = xor_cse_2608 ^ xor_cse_106 ^ xor_cse_286 ^ xor_cse_2855
      ^ Encrypt_Top_sbox_2_and_574 ^ state_1_1_63_32_lpi_4_24 ^ state_2_2_1_lpi_6;
  assign state_xor_808_nl = xor_cse_217 ^ xor_cse_218 ^ xor_cse_183 ^ xor_cse_285;
  assign state_xor_809_nl = xor_cse_1845 ^ xor_cse_1925 ^ (key1[25]) ^ xor_cse_389
      ^ xor_cse_1901;
  assign state_xor_810_nl = state_1_1_63_32_lpi_4_25 ^ state_2_3_1_lpi_4 ^ xor_cse_2610
      ^ xor_cse_293;
  assign state_xor_811_nl = state_1_1_63_32_lpi_4_25 ^ state_2_3_1_lpi_6 ^ xor_cse_2610
      ^ xor_cse_293;
  assign state_xor_812_nl = state_1_1_63_32_lpi_4_3 ^ xor_cse_228 ^ xor_cse_229 ^
      xor_cse_293;
  assign state_xor_813_nl = xor_cse_1868 ^ xor_cse_1919 ^ (key1[26]) ^ xor_cse_405
      ^ xor_cse_1913;
  assign state_xor_814_nl = state_1_1_63_32_lpi_4_26 ^ state_2_4_1_lpi_4 ^ xor_cse_2612
      ^ xor_cse_302;
  assign state_xor_815_nl = state_1_1_63_32_lpi_4_26 ^ state_2_4_1_lpi_6 ^ xor_cse_2612
      ^ xor_cse_302;
  assign state_xor_816_nl = state_1_1_63_32_lpi_4_30 ^ xor_cse_238 ^ xor_cse_239
      ^ xor_cse_302;
  assign state_xor_817_nl = xor_cse_1886 ^ xor_cse_1910 ^ (key1[27]) ^ xor_cse_417
      ^ xor_cse_1907;
  assign state_xor_818_nl = state_1_1_63_32_lpi_4_27 ^ state_2_5_1_lpi_4 ^ xor_cse_2618
      ^ xor_cse_311;
  assign state_xor_819_nl = state_1_1_63_32_lpi_4_27 ^ state_2_5_1_lpi_6 ^ xor_cse_2618
      ^ xor_cse_311;
  assign state_xor_820_nl = state_1_1_63_32_lpi_4_31 ^ xor_cse_248 ^ xor_cse_249
      ^ xor_cse_311;
  assign state_xor_821_nl = xor_cse_1895 ^ xor_cse_1898 ^ (key1[28]) ^ xor_cse_430
      ^ xor_cse_1892;
  assign state_xor_822_nl = state_1_1_63_32_lpi_4_28 ^ state_2_6_1_lpi_4 ^ xor_cse_2620
      ^ xor_cse_320;
  assign state_xor_823_nl = state_1_1_63_32_lpi_4_28 ^ state_2_6_1_lpi_6 ^ xor_cse_2620
      ^ xor_cse_320;
  assign state_xor_824_nl = state_1_1_63_32_lpi_4_4 ^ xor_cse_258 ^ xor_cse_260 ^
      xor_cse_320;
  assign state_xor_825_nl = xor_cse_1877 ^ xor_cse_1880 ^ (key1[29]) ^ xor_cse_444
      ^ xor_cse_1874;
  assign state_xor_826_nl = xor_cse_329 ^ (ROM_1i4_1o8_f17815f9d5076718618be5590cdd11c42e_1[7])
      ^ xor_cse_331 ^ state_1_1_63_32_lpi_4_29 ^ Encrypt_Top_sbox_2_and_576 ^ Encrypt_Top_sbox_2_and_578
      ^ state_2_7_1_lpi_4;
  assign state_xor_827_nl = state_1_1_63_32_lpi_4_29 ^ xor_cse_331 ^ xor_cse_2625
      ^ xor_cse_329;
  assign state_xor_828_nl = state_1_1_63_32_lpi_4_5 ^ xor_cse_270 ^ xor_cse_331 ^
      xor_cse_329;
  assign state_xor_667_nl = (key4[0]) ^ xor_cse_1735 ^ xor_cse_1736 ^ xor_cse_1737;
  assign state_xor_668_nl = xor_cse_148 ^ xor_cse_56 ^ xor_cse_2626 ^ state_4_4_0_lpi_3
      ^ state_4_4_7_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1;
  assign state_xor_670_nl = (key4[1]) ^ xor_cse_1742 ^ xor_cse_1743 ^ xor_cse_1744;
  assign state_xor_671_nl = xor_cse_70 ^ xor_cse_159 ^ xor_cse_2629 ^ state_4_4_1_lpi_3
      ^ state_4_4_8_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_42_sva_1;
  assign state_xor_673_nl = (key4[2]) ^ xor_cse_1749 ^ xor_cse_1750 ^ xor_cse_1751;
  assign state_xor_674_nl = xor_cse_84 ^ xor_cse_170 ^ xor_cse_151 ^ state_4_4_2_lpi_3
      ^ state_4_4_9_lpi_3 ^ state_4_4_43_lpi_3;
  assign state_xor_675_nl = (key4[3]) ^ xor_cse_1755 ^ xor_cse_1756 ^ xor_cse_1757;
  assign state_xor_676_nl = xor_cse_570 ^ xor_cse_569 ^ Encrypt_Top_sbox_1_and_cse_44_sva_1
      ^ state_3_44_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1 ^ state_1_1_63_32_lpi_4_12;
  assign state_xor_677_nl = (key4[4]) ^ xor_cse_1748 ^ xor_cse_1761 ^ xor_cse_1762;
  assign state_xor_678_nl = xor_cse_111 ^ xor_cse_168 ^ xor_cse_594 ^ state_4_4_4_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1 ^ state_4_4_45_lpi_3;
  assign state_xor_679_nl = (key4[5]) ^ xor_cse_1741 ^ xor_cse_1766 ^ xor_cse_1767;
  assign state_xor_680_nl = xor_cse_124 ^ xor_cse_181 ^ xor_cse_603 ^ xor_cse_605;
  assign state_xor_681_nl = (key4[6]) ^ xor_cse_1734 ^ xor_cse_1771 ^ xor_cse_1772;
  assign state_xor_682_nl = xor_cse_136 ^ xor_cse_192 ^ xor_cse_609 ^ state_4_4_6_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1 ^ state_4_4_47_lpi_3;
  assign state_xor_683_nl = (key4[7]) ^ xor_cse_1735 ^ xor_cse_1776 ^ xor_cse_1777;
  assign state_xor_684_nl = xor_cse_148 ^ xor_cse_201 ^ xor_cse_618 ^ state_4_4_7_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1 ^ state_4_4_48_lpi_3;
  assign state_xor_690_nl = xor_cse_1855 ^ xor_cse_1946 ^ xor_cse_401 ^ (key2[15])
      ^ xor_cse_1996 ^ xor_cse_1997 ^ state_4_3_63_32_sva_0;
  assign state_xor_691_nl = xor_cse_1357 ^ xor_cse_2641 ^ xor_cse_231 ^ xor_cse_1360;
  assign state_xor_692_nl = (key2[16]) ^ xor_cse_1835 ^ xor_cse_1955 ^ xor_cse_2001;
  assign state_xor_693_nl = xor_cse_2104 ^ xor_cse_242 ^ xor_cse_25 ^ xor_cse_2106
      ^ Encrypt_Top_sbox_2_and_758 ^ state_1_1_63_32_lpi_4_1;
  assign state_xor_694_nl = xor_cse_1963 ^ xor_cse_2008 ^ xor_cse_933 ^ (key2[17])
      ^ xor_cse_1853 ^ xor_cse_1854 ^ state_4_3_31_0_sva_17;
  assign state_xor_695_nl = xor_cse_2126 ^ xor_cse_1317 ^ xor_cse_252 ^ Encrypt_Top_sbox_2_and_658
      ^ state_4_4_17_lpi_3 ^ state_1_1_63_32_lpi_4_2;
  assign state_xor_696_nl = xor_cse_1871 ^ xor_cse_1970 ^ xor_cse_446 ^ (key2[18])
      ^ xor_cse_2018 ^ xor_cse_2019 ^ state_4_3_63_32_sva_3;
  assign state_xor_697_nl = xor_cse_1324 ^ xor_cse_2252 ^ xor_cse_263 ^ Encrypt_Top_sbox_2_and_666
      ^ state_4_4_18_lpi_3 ^ state_1_1_63_32_lpi_4_3;
  assign state_xor_698_nl = (key2[19]) ^ xor_cse_1889 ^ xor_cse_1976 ^ xor_cse_2025;
  assign state_xor_699_nl = xor_cse_2264 ^ xor_cse_2265 ^ xor_cse_369 ^ Encrypt_Top_sbox_2_and_754
      ^ state_4_4_29_lpi_3 ^ state_1_1_63_32_lpi_4_4;
  assign state_xor_700_nl = (key2[20]) ^ xor_cse_1904 ^ xor_cse_1982 ^ xor_cse_2033;
  assign state_xor_701_nl = xor_cse_1341 ^ xor_cse_2286 ^ xor_cse_282 ^ Encrypt_Top_sbox_2_and_682
      ^ state_4_4_20_lpi_3 ^ state_1_1_63_32_lpi_4_5;
  assign state_xor_702_nl = xor_cse_1916 ^ xor_cse_1988 ^ xor_cse_859 ^ (key2[21])
      ^ xor_cse_2041 ^ xor_cse_2042 ^ state_4_3_63_32_sva_6;
  assign state_xor_703_nl = xor_cse_1351 ^ xor_cse_1325 ^ xor_cse_92 ^ Encrypt_Top_sbox_2_and_716
      ^ Encrypt_Top_sbox_2_and_718 ^ state_1_1_63_32_lpi_4_6;
  assign state_xor_704_nl = xor_cse_1922 ^ xor_cse_2047 ^ xor_cse_401 ^ (key2[22])
      ^ xor_cse_1996 ^ xor_cse_1997 ^ state_4_3_63_32_sva_0;
  assign state_xor_705_nl = xor_cse_1332 ^ xor_cse_2641 ^ xor_cse_107 ^ Encrypt_Top_sbox_2_and_708
      ^ Encrypt_Top_sbox_2_and_710 ^ state_1_1_63_32_lpi_4_7;
  assign state_xor_706_nl = xor_cse_1928 ^ xor_cse_2001 ^ xor_cse_878 ^ (key2[23])
      ^ xor_cse_2054 ^ xor_cse_2055 ^ state_4_3_63_32_sva_8;
  assign state_xor_707_nl = xor_cse_2315 ^ xor_cse_2316 ^ xor_cse_120 ^ state_1_1_63_32_lpi_4_1
      ^ Encrypt_Top_sbox_2_and_702 ^ state_1_1_63_32_lpi_4_8;
  assign state_xor_708_nl = xor_cse_1936 ^ xor_cse_2008 ^ xor_cse_888 ^ (key2[24])
      ^ xor_cse_2045 ^ xor_cse_2046 ^ state_4_3_63_32_sva_9;
  assign state_xor_709_nl = xor_cse_1350 ^ xor_cse_130 ^ xor_cse_38 ^ Encrypt_Top_sbox_2_and_748
      ^ Encrypt_Top_sbox_2_and_750 ^ state_1_1_63_32_lpi_4_2 ^ Encrypt_Top_sbox_2_and_692
      ^ Encrypt_Top_sbox_2_and_694 ^ state_1_1_63_32_lpi_4_9;
  assign state_xor_710_nl = xor_cse_1946 ^ xor_cse_2036 ^ xor_cse_446 ^ (key2[25])
      ^ xor_cse_2018 ^ xor_cse_2019 ^ state_4_3_63_32_sva_3;
  assign state_xor_711_nl = xor_cse_1357 ^ xor_cse_8 ^ xor_cse_52 ^ Encrypt_Top_sbox_2_and_740
      ^ Encrypt_Top_sbox_2_and_742 ^ state_1_1_63_32_lpi_4_3 ^ Encrypt_Top_sbox_2_and_684
      ^ Encrypt_Top_sbox_2_and_686 ^ state_1_1_63_32_lpi_4_10;
  assign state_xor_712_nl = xor_cse_1955 ^ xor_cse_2025 ^ xor_cse_910 ^ (key2[26])
      ^ xor_cse_2030 ^ xor_cse_2032 ^ state_4_3_63_32_sva_11;
  assign state_xor_713_nl = xor_cse_2104 ^ xor_cse_22 ^ xor_cse_66 ^ Encrypt_Top_sbox_2_and_732
      ^ Encrypt_Top_sbox_2_and_734 ^ state_1_1_63_32_lpi_4_4 ^ Encrypt_Top_sbox_2_and_676
      ^ Encrypt_Top_sbox_2_and_678 ^ state_1_1_63_32_lpi_4_11;
  assign state_xor_714_nl = xor_cse_1963 ^ xor_cse_2033 ^ xor_cse_924 ^ (key2[27])
      ^ xor_cse_2022 ^ xor_cse_2024 ^ state_4_3_63_32_sva_12;
  assign state_xor_715_nl = xor_cse_1317 ^ xor_cse_2688 ^ xor_cse_80 ^ Encrypt_Top_sbox_2_and_724
      ^ Encrypt_Top_sbox_2_and_726 ^ state_1_1_63_32_lpi_4_5;
  assign state_xor_716_nl = xor_cse_1970 ^ xor_cse_2013 ^ xor_cse_859 ^ (key2[28])
      ^ xor_cse_2041 ^ xor_cse_2042 ^ state_4_3_63_32_sva_6;
  assign state_xor_717_nl = xor_cse_1324 ^ xor_cse_49 ^ xor_cse_92 ^ Encrypt_Top_sbox_2_and_716
      ^ Encrypt_Top_sbox_2_and_718 ^ state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_2_and_660
      ^ Encrypt_Top_sbox_2_and_662 ^ state_1_1_63_32_lpi_4_13;
  assign state_xor_718_nl = xor_cse_1976 ^ xor_cse_2047 ^ xor_cse_948 ^ (key2[29])
      ^ xor_cse_2006 ^ xor_cse_2007 ^ state_4_3_63_32_sva_14;
  assign state_xor_719_nl = xor_cse_2367 ^ xor_cse_63 ^ xor_cse_369 ^ Encrypt_Top_sbox_2_and_754
      ^ state_4_4_29_lpi_3 ^ state_1_1_63_32_lpi_4_7 ^ Encrypt_Top_sbox_2_and_652
      ^ Encrypt_Top_sbox_2_and_654 ^ state_1_1_63_32_lpi_4_14;
  assign state_xor_720_nl = xor_cse_1982 ^ xor_cse_1998 ^ xor_cse_878 ^ (key2[30])
      ^ xor_cse_2054 ^ xor_cse_2055 ^ state_4_3_63_32_sva_8;
  assign state_xor_721_nl = xor_cse_1341 ^ xor_cse_2379 ^ xor_cse_77 ^ state_1_1_63_32_lpi_4_8
      ^ Encrypt_Top_sbox_2_and_646 ^ state_1_1_63_32_lpi_4_15;
  assign state_xor_722_nl = xor_cse_1988 ^ xor_cse_1991 ^ xor_cse_888 ^ (key2[31])
      ^ xor_cse_2045 ^ xor_cse_2046 ^ state_4_3_63_32_sva_9;
  assign state_xor_723_nl = xor_cse_2707 ^ xor_cse_1351 ^ xor_cse_130 ^ Encrypt_Top_sbox_2_and_692
      ^ Encrypt_Top_sbox_2_and_694 ^ state_1_1_63_32_lpi_4_9;
  assign state_xor_724_nl = xor_cse_2036 ^ xor_cse_1985 ^ xor_cse_401 ^ xor_cse_1996
      ^ xor_cse_1997 ^ state_4_3_63_32_sva_0 ^ (key1[0]);
  assign state_xor_725_nl = xor_cse_7 ^ xor_cse_10 ^ xor_cse_11 ^ Encrypt_Top_sbox_2_and_764
      ^ state_1_1_63_32_lpi_4_0 ^ state_1_1_63_32_lpi_4_10 ^ Encrypt_Top_sbox_2_and_628
      ^ Encrypt_Top_sbox_2_and_630 ^ state_1_1_63_32_lpi_4_17;
  assign state_xor_726_nl = xor_cse_7 ^ xor_cse_10 ^ xor_cse_11 ^ xor_cse_12 ^ state_1_1_31_0_lpi_4_8
      ^ state_1_1_63_32_lpi_4_16;
  assign state_xor_727_nl = xor_cse_1979 ^ xor_cse_2001 ^ xor_cse_910 ^ xor_cse_2030
      ^ xor_cse_2032 ^ state_4_3_63_32_sva_11 ^ (key1[1]);
  assign state_xor_728_nl = xor_cse_21 ^ xor_cse_24 ^ xor_cse_25 ^ Encrypt_Top_sbox_2_and_620
      ^ Encrypt_Top_sbox_2_and_756 ^ state_1_1_63_32_lpi_4_1 ^ state_1_1_63_32_lpi_4_11
      ^ Encrypt_Top_sbox_2_and_622 ^ state_1_1_63_32_lpi_4_18;
  assign state_xor_729_nl = xor_cse_21 ^ xor_cse_24 ^ xor_cse_25 ^ xor_cse_26 ^ state_1_1_31_0_lpi_4_9
      ^ state_1_1_63_32_lpi_4_17;
  assign state_xor_730_nl = xor_cse_1973 ^ xor_cse_2008 ^ xor_cse_924 ^ xor_cse_2022
      ^ xor_cse_2024 ^ state_4_3_63_32_sva_12 ^ (key1[2]);
  assign state_xor_731_nl = xor_cse_2688 ^ xor_cse_37 ^ xor_cse_38 ^ Encrypt_Top_sbox_2_and_612
      ^ Encrypt_Top_sbox_2_and_614 ^ Encrypt_Top_sbox_2_and_748 ^ Encrypt_Top_sbox_2_and_750
      ^ state_1_1_63_32_lpi_4_2 ^ state_1_1_63_32_lpi_4_19;
  assign state_xor_732_nl = xor_cse_34 ^ xor_cse_37 ^ xor_cse_38 ^ xor_cse_39 ^ Encrypt_Top_sbox_2_and_750
      ^ state_1_1_63_32_lpi_4_0;
  assign state_xor_733_nl = xor_cse_1966 ^ xor_cse_2013 ^ xor_cse_446 ^ xor_cse_2018
      ^ xor_cse_2019 ^ state_4_3_63_32_sva_3 ^ (key1[3]);
  assign state_xor_734_nl = xor_cse_48 ^ xor_cse_51 ^ xor_cse_52 ^ Encrypt_Top_sbox_2_and_740
      ^ state_1_1_63_32_lpi_4_3 ^ state_1_1_63_32_lpi_4_13 ^ Encrypt_Top_sbox_2_and_604
      ^ Encrypt_Top_sbox_2_and_606 ^ state_1_1_63_32_lpi_4_20;
  assign state_xor_735_nl = xor_cse_48 ^ xor_cse_51 ^ xor_cse_52 ^ xor_cse_53 ^ state_1_1_63_32_lpi_4_1
      ^ state_1_1_63_32_lpi_4_19;
  assign state_xor_736_nl = xor_cse_1960 ^ xor_cse_2025 ^ xor_cse_948 ^ xor_cse_2006
      ^ xor_cse_2007 ^ state_4_3_63_32_sva_14 ^ (key1[4]);
  assign state_xor_737_nl = xor_cse_62 ^ xor_cse_65 ^ xor_cse_66 ^ Encrypt_Top_sbox_2_and_732
      ^ state_1_1_63_32_lpi_4_4 ^ state_1_1_63_32_lpi_4_14 ^ Encrypt_Top_sbox_2_and_596
      ^ Encrypt_Top_sbox_2_and_598 ^ state_1_1_63_32_lpi_4_21;
  assign state_xor_738_nl = xor_cse_62 ^ xor_cse_65 ^ xor_cse_66 ^ xor_cse_67 ^ state_1_1_63_32_lpi_4_10
      ^ state_1_1_63_32_lpi_4_2;
  assign state_xor_739_nl = (key1[5]) ^ xor_cse_1951 ^ xor_cse_1998 ^ xor_cse_2033;
  assign state_xor_740_nl = xor_cse_76 ^ xor_cse_79 ^ xor_cse_80 ^ Encrypt_Top_sbox_2_and_588
      ^ Encrypt_Top_sbox_2_and_590 ^ Encrypt_Top_sbox_2_and_724 ^ state_1_1_63_32_lpi_4_5
      ^ state_1_1_63_32_lpi_4_15 ^ state_1_1_63_32_lpi_4_22;
  assign state_xor_741_nl = xor_cse_76 ^ xor_cse_79 ^ xor_cse_80 ^ xor_cse_81 ^ state_1_1_63_32_lpi_4_11
      ^ state_1_1_63_32_lpi_4_20;
  assign state_xor_742_nl = xor_cse_1941 ^ xor_cse_1991 ^ xor_cse_859 ^ xor_cse_2041
      ^ xor_cse_2042 ^ state_4_3_63_32_sva_6 ^ (key1[6]);
  assign state_xor_743_nl = xor_cse_2707 ^ xor_cse_91 ^ xor_cse_92 ^ Encrypt_Top_sbox_2_and_716
      ^ Encrypt_Top_sbox_2_and_718 ^ state_1_1_63_32_lpi_4_6 ^ Encrypt_Top_sbox_2_and_580
      ^ Encrypt_Top_sbox_2_and_582 ^ state_1_1_63_32_lpi_4_23;
  assign state_xor_744_nl = xor_cse_90 ^ xor_cse_94 ^ xor_cse_95 ^ xor_cse_2387;
  assign state_xor_745_nl = (key1[7]) ^ xor_cse_1931 ^ xor_cse_1985 ^ xor_cse_2047;
  assign state_xor_746_nl = xor_cse_104 ^ xor_cse_106 ^ xor_cse_107 ^ Encrypt_Top_sbox_2_and_708
      ^ state_1_1_63_32_lpi_4_7 ^ state_1_1_63_32_lpi_4_17 ^ Encrypt_Top_sbox_2_and_572
      ^ Encrypt_Top_sbox_2_and_574 ^ state_1_1_63_32_lpi_4_24;
  assign state_xor_747_nl = xor_cse_104 ^ xor_cse_106 ^ xor_cse_107 ^ xor_cse_108
      ^ state_1_1_63_32_lpi_4_13 ^ state_1_1_63_32_lpi_4_22;
  assign state_xor_748_nl = xor_cse_1925 ^ xor_cse_1979 ^ xor_cse_878 ^ xor_cse_2054
      ^ xor_cse_2055 ^ state_4_3_63_32_sva_8 ^ (key1[8]);
  assign state_xor_749_nl = xor_cse_117 ^ xor_cse_119 ^ xor_cse_120 ^ Encrypt_Top_sbox_2_and_700
      ^ Encrypt_Top_sbox_2_and_564 ^ Encrypt_Top_sbox_2_and_566 ^ state_1_1_63_32_lpi_4_8
      ^ state_1_1_63_32_lpi_4_18 ^ state_1_1_63_32_lpi_4_25;
  assign state_xor_750_nl = xor_cse_117 ^ xor_cse_119 ^ xor_cse_120 ^ xor_cse_121
      ^ state_1_1_63_32_lpi_4_14 ^ state_1_1_63_32_lpi_4_23;
  assign state_xor_751_nl = xor_cse_1919 ^ xor_cse_1973 ^ xor_cse_888 ^ xor_cse_2045
      ^ xor_cse_2046 ^ state_4_3_63_32_sva_9 ^ (key1[9]);
  assign state_xor_752_nl = xor_cse_2771 ^ xor_cse_129 ^ xor_cse_37 ^ Encrypt_Top_sbox_2_and_692
      ^ state_1_1_63_32_lpi_4_9 ^ state_1_1_63_32_lpi_4_19;
  assign state_xor_753_nl = xor_cse_129 ^ xor_cse_132 ^ xor_cse_37 ^ xor_cse_133
      ^ state_1_1_63_32_lpi_4_15 ^ state_1_1_63_32_lpi_4_24;
  assign state_xor_754_nl = (key1[10]) ^ xor_cse_1910 ^ xor_cse_1966 ^ xor_cse_2036;
  assign state_xor_755_nl = xor_cse_143 ^ xor_cse_142 ^ Encrypt_Top_sbox_2_and_548
      ^ Encrypt_Top_sbox_2_and_684 ^ Encrypt_Top_sbox_2_and_686 ^ state_1_1_63_32_lpi_4_10
      ^ Encrypt_Top_sbox_2_and_604 ^ state_1_1_63_32_lpi_4_20 ^ Encrypt_Top_sbox_2_and_550
      ^ state_1_1_63_32_lpi_4_27;
  assign state_xor_756_nl = state_1_1_63_32_lpi_4_25 ^ xor_cse_145 ^ xor_cse_141
      ^ xor_cse_143;
  assign state_xor_757_nl = xor_cse_1960 ^ xor_cse_910 ^ xor_cse_1528 ^ xor_cse_2029
      ^ xor_cse_2032 ^ state_4_3_63_32_sva_11 ^ (key1[11]);
  assign state_xor_758_nl = state_1_1_63_32_lpi_4_28 ^ xor_cse_154 ^ xor_cse_65 ^
      xor_cse_22 ^ Encrypt_Top_sbox_2_and_540 ^ Encrypt_Top_sbox_2_and_542 ^ Encrypt_Top_sbox_2_and_676
      ^ Encrypt_Top_sbox_2_and_678 ^ state_1_1_63_32_lpi_4_11 ^ Encrypt_Top_sbox_2_and_596
      ^ Encrypt_Top_sbox_2_and_598 ^ state_1_1_63_32_lpi_4_21;
  assign state_xor_759_nl = xor_cse_153 ^ xor_cse_65 ^ xor_cse_22 ^ xor_cse_156 ^
      Encrypt_Top_sbox_2_and_598 ^ state_1_1_63_32_lpi_4_26;
  assign state_xor_760_nl = xor_cse_1951 ^ xor_cse_924 ^ xor_cse_1375 ^ xor_cse_2021
      ^ xor_cse_2024 ^ state_4_3_63_32_sva_12 ^ (key1[12]);
  assign state_xor_761_nl = xor_cse_163 ^ xor_cse_2688 ^ xor_cse_79 ^ state_1_1_63_32_lpi_4_22
      ^ Encrypt_Top_sbox_2_and_532 ^ state_1_1_63_32_lpi_4_29;
  assign state_xor_762_nl = xor_cse_34 ^ xor_cse_163 ^ xor_cse_79 ^ state_1_1_63_32_lpi_4_27
      ^ Encrypt_Top_sbox_2_and_532 ^ state_1_1_63_32_lpi_4_5;
  assign state_xor_763_nl = (key1[13]) ^ xor_cse_1941 ^ xor_cse_2013 ^ xor_cse_1969;
  assign state_xor_764_nl = xor_cse_2791 ^ xor_cse_91 ^ xor_cse_49 ^ Encrypt_Top_sbox_2_and_524
      ^ Encrypt_Top_sbox_2_and_660 ^ Encrypt_Top_sbox_2_and_662 ^ state_1_1_63_32_lpi_4_13
      ^ Encrypt_Top_sbox_2_and_580 ^ Encrypt_Top_sbox_2_and_582 ^ state_1_1_63_32_lpi_4_23;
  assign state_xor_765_nl = xor_cse_172 ^ xor_cse_174 ^ xor_cse_49 ^ xor_cse_175
      ^ Encrypt_Top_sbox_2_and_662 ^ state_1_1_63_32_lpi_4_19;
  assign state_xor_766_nl = xor_cse_1838 ^ xor_cse_1931 ^ xor_cse_948 ^ xor_cse_2006
      ^ xor_cse_2007 ^ state_4_3_63_32_sva_14 ^ (key1[14]);
  assign state_xor_767_nl = xor_cse_2799 ^ xor_cse_106 ^ xor_cse_63 ^ Encrypt_Top_sbox_2_and_516
      ^ Encrypt_Top_sbox_2_and_652 ^ Encrypt_Top_sbox_2_and_654 ^ state_1_1_63_32_lpi_4_14
      ^ Encrypt_Top_sbox_2_and_572 ^ Encrypt_Top_sbox_2_and_574 ^ state_1_1_63_32_lpi_4_24;
  assign state_xor_768_nl = xor_cse_183 ^ xor_cse_185 ^ xor_cse_63 ^ xor_cse_186
      ^ xor_cse_2370;
  assign state_xor_829_nl = xor_cse_1855 ^ xor_cse_1162 ^ xor_cse_1400 ^ xor_cse_1859
      ^ xor_cse_1864 ^ state_4_3_31_0_sva_8 ^ (key1[30]);
  assign state_xor_830_nl = xor_cse_231 ^ xor_cse_339 ^ xor_cse_2791 ^ xor_cse_2868;
  assign state_xor_831_nl = xor_cse_277 ^ xor_cse_174 ^ xor_cse_231 ^ xor_cse_339
      ^ Encrypt_Top_sbox_2_and_526 ^ state_1_1_63_32_lpi_4_6;
  assign state_xor_832_nl = xor_cse_1835 ^ xor_cse_1838 ^ xor_cse_1172 ^ xor_cse_1843
      ^ xor_cse_1844 ^ state_4_3_31_0_sva_9 ^ (key1[31]);
  assign state_xor_833_nl = xor_cse_2799 ^ xor_cse_286 ^ xor_cse_242 ^ xor_cse_347
      ^ Encrypt_Top_sbox_2_and_592 ^ Encrypt_Top_sbox_2_and_594 ^ state_1_1_31_0_lpi_4_9;
  assign state_xor_834_nl = xor_cse_285 ^ xor_cse_185 ^ xor_cse_242 ^ xor_cse_347
      ^ Encrypt_Top_sbox_2_and_518 ^ state_1_1_63_32_lpi_4_7;
  assign state_xor_835_nl = xor_cse_1871 ^ xor_cse_1946 ^ xor_cse_1162 ^ (key2[8])
      ^ xor_cse_1862 ^ xor_cse_1864 ^ state_4_3_31_0_sva_8;
  assign state_xor_836_nl = xor_cse_1357 ^ xor_cse_2868 ^ xor_cse_263 ^ xor_cse_2421;
  assign state_xor_837_nl = xor_cse_1889 ^ xor_cse_1955 ^ xor_cse_1172 ^ (key2[9])
      ^ xor_cse_1843 ^ xor_cse_1844 ^ state_4_3_31_0_sva_9;
  assign state_xor_838_nl = xor_cse_2104 ^ xor_cse_286 ^ xor_cse_274 ^ Encrypt_Top_sbox_2_and_592
      ^ Encrypt_Top_sbox_2_and_594 ^ state_1_1_31_0_lpi_4_9 ^ Encrypt_Top_sbox_2_and_672
      ^ Encrypt_Top_sbox_2_and_674 ^ state_4_4_19_lpi_3;
  assign state_xor_839_nl = xor_cse_861 ^ xor_cse_1789 ^ xor_cse_1790 ^ (key4[10])
      ^ state_4_3_31_0_sva_10 ^ Encrypt_Top_sbox_and_2_cse_17_sva_1 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1;
  assign state_xor_840_nl = xor_cse_1 ^ xor_cse_479 ^ xor_cse_569 ^ xor_cse_2887;
  assign state_xor_842_nl = (key4[11]) ^ xor_cse_868 ^ xor_cse_1792 ^ xor_cse_1794;
  assign state_xor_843_nl = xor_cse_15 ^ xor_cse_594 ^ xor_cse_491 ^ xor_cse_2889;
  assign state_xor_845_nl = (key4[12]) ^ xor_cse_880 ^ xor_cse_1787 ^ xor_cse_1796;
  assign state_xor_846_nl = xor_cse_29 ^ xor_cse_603 ^ xor_cse_498 ^ xor_cse_2891;
  assign state_xor_848_nl = (key4[13]) ^ xor_cse_890 ^ xor_cse_1783 ^ xor_cse_1798;
  assign state_xor_849_nl = xor_cse_44 ^ xor_cse_609 ^ xor_cse_514 ^ xor_cse_2893;
  assign state_xor_851_nl = (key4[14]) ^ xor_cse_900 ^ xor_cse_1778 ^ xor_cse_1800;
  assign state_xor_852_nl = xor_cse_57 ^ xor_cse_618 ^ xor_cse_520 ^ xor_cse_2895;
  assign state_xor_854_nl = (key4[15]) ^ xor_cse_1773 ^ xor_cse_912 ^ xor_cse_1802;
  assign state_xor_855_nl = xor_cse_73 ^ xor_cse_673 ^ xor_cse_528 ^ xor_cse_2897;
  assign state_xor_857_nl = (key4[16]) ^ xor_cse_926 ^ xor_cse_1768 ^ xor_cse_1804;
  assign state_xor_858_nl = xor_cse_85 ^ xor_cse_468 ^ xor_cse_469 ^ xor_cse_471;
  assign state_xor_859_nl = xor_cse_415 ^ xor_cse_1790 ^ xor_cse_1763 ^ (key4[17])
      ^ Encrypt_Top_sbox_and_2_cse_17_sva_1 ^ state_4_3_31_0_sva_24 ^ Encrypt_Top_sbox_and_2_cse_58_sva_1;
  assign state_xor_860_nl = xor_cse_100 ^ xor_cse_479 ^ xor_cse_481 ^ xor_cse_482;
  assign state_xor_861_nl = xor_cse_428 ^ xor_cse_951 ^ xor_cse_1758 ^ (key4[18])
      ^ state_4_3_31_0_sva_18 ^ state_4_3_31_0_sva_25 ^ Encrypt_Top_sbox_and_2_cse_59_sva_1;
  assign state_xor_862_nl = xor_cse_490 ^ xor_cse_491 ^ xor_cse_2903 ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1;
  assign state_xor_863_nl = xor_cse_1078 ^ xor_cse_350 ^ xor_cse_448 ^ (key4[19])
      ^ state_4_3_31_0_sva_19 ^ state_4_3_31_0_sva_26 ^ state_4_3_63_32_sva_28;
  assign state_xor_864_nl = xor_cse_498 ^ xor_cse_500 ^ xor_cse_2906 ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_26_sva_1 ^ state_3_60_lpi_3;
  assign state_xor_865_nl = xor_cse_1087 ^ xor_cse_362 ^ xor_cse_1031 ^ (key4[20])
      ^ state_4_3_31_0_sva_20 ^ state_4_3_31_0_sva_27 ^ state_4_3_63_32_sva_29;
  assign state_xor_866_nl = xor_cse_514 ^ xor_cse_516 ^ xor_cse_2909 ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1
      ^ state_1_1_31_0_lpi_4_27 ^ state_3_61_lpi_3;
  assign state_xor_867_nl = xor_cse_1097 ^ xor_cse_354 ^ xor_cse_375 ^ (key4[21])
      ^ state_4_3_31_0_sva_21 ^ state_4_3_31_0_sva_28 ^ state_4_3_63_32_sva_30;
  assign state_xor_868_nl = xor_cse_520 ^ xor_cse_522 ^ xor_cse_2912 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1
      ^ Encrypt_Top_sbox_2_and_2_cse_28_sva_1 ^ state_1_1_63_32_lpi_4_30;
  assign state_xor_869_nl = xor_cse_366 ^ xor_cse_387 ^ xor_cse_1732 ^ (key4[22])
      ^ state_4_3_31_0_sva_22 ^ state_4_3_31_0_sva_29 ^ Encrypt_Top_sbox_and_2_cse_63_sva_1;
  assign state_xor_870_nl = xor_cse_42 ^ xor_cse_526 ^ xor_cse_528 ^ xor_cse_529;
  assign state_xor_873_nl = xor_cse_1752 ^ xor_cse_428 ^ xor_cse_1780 ^ (key4[25])
      ^ state_4_3_31_0_sva_25 ^ Encrypt_Top_sbox_and_2_cse_32_sva_1 ^ Encrypt_Top_sbox_and_2_cse_2_sva_1;
  assign state_xor_874_nl = xor_cse_84 ^ xor_cse_4 ^ xor_cse_490 ^ xor_cse_542;
  assign state_xor_875_nl = xor_cse_1755 ^ xor_cse_448 ^ xor_cse_1775 ^ (key4[26])
      ^ state_4_3_31_0_sva_26 ^ Encrypt_Top_sbox_and_2_cse_33_sva_1 ^ Encrypt_Top_sbox_and_2_cse_3_sva_1;
  assign state_xor_876_nl = xor_cse_102 ^ xor_cse_18 ^ xor_cse_500 ^ xor_cse_547;
  assign state_xor_877_nl = xor_cse_1748 ^ xor_cse_1031 ^ xor_cse_1770 ^ (key4[27])
      ^ state_4_3_31_0_sva_27 ^ Encrypt_Top_sbox_and_2_cse_34_sva_1 ^ Encrypt_Top_sbox_and_2_cse_4_sva_1;
  assign state_xor_878_nl = xor_cse_111 ^ xor_cse_30 ^ xor_cse_516 ^ xor_cse_552;
  assign state_xor_879_nl = xor_cse_1741 ^ xor_cse_354 ^ xor_cse_1765 ^ (key4[28])
      ^ state_4_3_31_0_sva_28 ^ Encrypt_Top_sbox_and_2_cse_35_sva_1 ^ Encrypt_Top_sbox_and_2_cse_5_sva_1;
  assign state_xor_880_nl = xor_cse_124 ^ xor_cse_46 ^ xor_cse_522 ^ xor_cse_557;
  assign state_xor_881_nl = xor_cse_1734 ^ xor_cse_366 ^ xor_cse_1760 ^ (key4[29])
      ^ state_4_3_31_0_sva_29 ^ Encrypt_Top_sbox_and_2_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_6_sva_1;
  assign state_xor_882_nl = xor_cse_59 ^ xor_cse_526 ^ xor_cse_562;
  assign state_xor_883_nl = xor_cse_1735 ^ xor_cse_379 ^ xor_cse_1753 ^ (key4[30])
      ^ state_4_3_31_0_sva_30 ^ Encrypt_Top_sbox_and_2_cse_37_sva_1 ^ Encrypt_Top_sbox_and_2_cse_7_sva_1;
  assign state_xor_884_nl = xor_cse_577 ^ xor_cse_74 ^ state_3_30_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_30_sva_1
      ^ state_1_1_31_0_lpi_4_30 ^ state_4_4_37_lpi_3;
  assign state_xor_885_nl = xor_cse_390 ^ xor_cse_1746 ^ xor_cse_1743 ^ (key4[31])
      ^ state_4_3_31_0_sva_31 ^ Encrypt_Top_sbox_and_2_cse_38_sva_1 ^ Encrypt_Top_sbox_and_2_cse_8_sva_1;
  assign state_xor_886_nl = xor_cse_159 ^ xor_cse_87 ^ xor_cse_536 ^ xor_cse_589;
  assign state_xor_887_nl = xor_cse_1739 ^ xor_cse_1780 ^ xor_cse_1750 ^ (key3[0])
      ^ Encrypt_Top_sbox_and_2_cse_32_sva_1 ^ Encrypt_Top_sbox_and_2_cse_39_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_9_sva_1;
  assign state_xor_888_nl = xor_cse_170 ^ xor_cse_98 ^ xor_cse_4 ^ state_4_4_32_lpi_3
      ^ state_4_4_39_lpi_3 ^ state_4_4_9_lpi_3;
  assign state_xor_889_nl = xor_cse_1731 ^ xor_cse_861 ^ xor_cse_1775 ^ (key3[1])
      ^ Encrypt_Top_sbox_and_2_cse_33_sva_1 ^ Encrypt_Top_sbox_and_2_cse_40_sva_1
      ^ state_4_3_31_0_sva_10;
  assign state_xor_890_nl = xor_cse_113 ^ xor_cse_18 ^ xor_cse_569 ^ xor_cse_636;
  assign state_xor_891_nl = xor_cse_1736 ^ xor_cse_868 ^ xor_cse_1770 ^ (key3[2])
      ^ Encrypt_Top_sbox_and_2_cse_34_sva_1 ^ Encrypt_Top_sbox_and_2_cse_41_sva_1
      ^ state_4_3_31_0_sva_11;
  assign state_xor_892_nl = xor_cse_30 ^ xor_cse_594 ^ xor_cse_2626 ^ state_4_4_34_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_11_sva_1;
  assign state_xor_893_nl = xor_cse_1742 ^ xor_cse_880 ^ xor_cse_1765 ^ (key3[3])
      ^ Encrypt_Top_sbox_and_2_cse_35_sva_1 ^ Encrypt_Top_sbox_and_2_cse_42_sva_1
      ^ state_4_3_31_0_sva_12;
  assign state_xor_894_nl = xor_cse_46 ^ xor_cse_603 ^ xor_cse_2629 ^ state_4_4_35_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_42_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_12_sva_1;
  assign state_xor_895_nl = xor_cse_1749 ^ xor_cse_890 ^ xor_cse_1760 ^ (key3[4])
      ^ Encrypt_Top_sbox_and_2_cse_36_sva_1 ^ Encrypt_Top_sbox_and_2_cse_43_sva_1
      ^ state_4_3_31_0_sva_13;
  assign state_xor_896_nl = xor_cse_151 ^ xor_cse_59 ^ xor_cse_609 ^ state_4_4_36_lpi_3
      ^ state_4_4_43_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_13_sva_1;
  assign state_xor_897_nl = xor_cse_1756 ^ xor_cse_900 ^ xor_cse_1753 ^ (key3[5])
      ^ Encrypt_Top_sbox_and_2_cse_37_sva_1 ^ Encrypt_Top_sbox_and_2_cse_44_sva_1
      ^ state_4_3_31_0_sva_14;
  assign state_xor_898_nl = xor_cse_74 ^ xor_cse_618 ^ state_4_4_37_lpi_3 ^ Encrypt_Top_sbox_1_and_cse_44_sva_1
      ^ state_4_4_44_lpi_3 ^ state_3_44_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1
      ^ state_1_1_63_32_lpi_4_12 ^ Encrypt_Top_sbox_2_and_2_cse_14_sva_1;
  assign state_xor_899_nl = xor_cse_1761 ^ xor_cse_912 ^ xor_cse_1746 ^ (key3[6])
      ^ Encrypt_Top_sbox_and_2_cse_38_sva_1 ^ Encrypt_Top_sbox_and_2_cse_45_sva_1
      ^ state_4_3_31_0_sva_15;
  assign state_xor_900_nl = xor_cse_168 ^ xor_cse_87 ^ xor_cse_673 ^ state_4_4_38_lpi_3
      ^ state_4_4_45_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_15_sva_1;
  assign state_xor_901_nl = xor_cse_1739 ^ xor_cse_926 ^ xor_cse_1766 ^ (key3[7])
      ^ Encrypt_Top_sbox_and_2_cse_39_sva_1 ^ Encrypt_Top_sbox_and_2_cse_46_sva_1
      ^ state_4_3_31_0_sva_16;
  assign state_xor_902_nl = xor_cse_98 ^ xor_cse_181 ^ xor_cse_469 ^ state_4_4_39_lpi_3
      ^ state_4_4_46_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1;
  assign state_xor_903_nl = xor_cse_1731 ^ xor_cse_1771 ^ xor_cse_1790 ^ (key3[8])
      ^ Encrypt_Top_sbox_and_2_cse_40_sva_1 ^ Encrypt_Top_sbox_and_2_cse_47_sva_1
      ^ Encrypt_Top_sbox_and_2_cse_17_sva_1;
  assign state_xor_904_nl = xor_cse_192 ^ xor_cse_113 ^ xor_cse_479 ^ state_4_4_40_lpi_3
      ^ state_4_4_47_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_17_sva_1;
  assign state_xor_905_nl = xor_cse_1736 ^ xor_cse_951 ^ xor_cse_1776 ^ (key3[9])
      ^ Encrypt_Top_sbox_and_2_cse_41_sva_1 ^ Encrypt_Top_sbox_and_2_cse_48_sva_1
      ^ state_4_3_31_0_sva_18;
  assign state_xor_906_nl = xor_cse_201 ^ xor_cse_491 ^ xor_cse_2626 ^ Encrypt_Top_sbox_2_and_2_cse_41_sva_1
      ^ state_4_4_48_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_18_sva_1;
  assign state_xor_907_nl = xor_cse_1742 ^ xor_cse_350 ^ xor_cse_1781 ^ (key3[10])
      ^ Encrypt_Top_sbox_and_2_cse_42_sva_1 ^ Encrypt_Top_sbox_and_2_cse_49_sva_1
      ^ state_4_3_31_0_sva_19;
  assign state_xor_908_nl = xor_cse_214 ^ xor_cse_498 ^ xor_cse_2629 ^ Encrypt_Top_sbox_2_and_2_cse_42_sva_1
      ^ state_4_4_49_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_19_sva_1;
  assign state_xor_909_nl = xor_cse_1749 ^ xor_cse_362 ^ xor_cse_1785 ^ (key3[11])
      ^ Encrypt_Top_sbox_and_2_cse_43_sva_1 ^ Encrypt_Top_sbox_and_2_cse_50_sva_1
      ^ state_4_3_31_0_sva_20;
  assign state_xor_910_nl = xor_cse_224 ^ xor_cse_151 ^ xor_cse_514 ^ state_4_4_43_lpi_3
      ^ state_4_4_50_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_20_sva_1;
  assign state_xor_911_nl = xor_cse_1756 ^ xor_cse_375 ^ xor_cse_1789 ^ (key3[12])
      ^ Encrypt_Top_sbox_and_2_cse_44_sva_1 ^ Encrypt_Top_sbox_and_2_cse_51_sva_1
      ^ state_4_3_31_0_sva_21;
  assign state_xor_912_nl = xor_cse_1 ^ xor_cse_520 ^ Encrypt_Top_sbox_1_and_cse_44_sva_1
      ^ state_4_4_44_lpi_3 ^ state_3_44_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_44_sva_1
      ^ state_1_1_63_32_lpi_4_12 ^ state_4_4_51_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_21_sva_1;
  assign state_xor_913_nl = xor_cse_1761 ^ xor_cse_387 ^ xor_cse_1792 ^ (key3[13])
      ^ Encrypt_Top_sbox_and_2_cse_45_sva_1 ^ Encrypt_Top_sbox_and_2_cse_52_sva_1
      ^ state_4_3_31_0_sva_22;
  assign state_xor_914_nl = xor_cse_15 ^ xor_cse_168 ^ xor_cse_528 ^ state_4_4_45_lpi_3
      ^ state_4_4_52_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_22_sva_1;
  assign state_xor_915_nl = xor_cse_403 ^ xor_cse_1766 ^ xor_cse_1787 ^ (key3[14])
      ^ Encrypt_Top_sbox_and_2_cse_46_sva_1 ^ Encrypt_Top_sbox_and_2_cse_53_sva_1
      ^ state_4_3_31_0_sva_23;
  assign state_xor_916_nl = xor_cse_29 ^ xor_cse_181 ^ xor_cse_468 ^ xor_cse_735;
  assign state_xor_917_nl = (key3[15]) ^ xor_cse_1771 ^ xor_cse_1783 ^ xor_cse_1803;
  assign state_xor_918_nl = xor_cse_44 ^ xor_cse_192 ^ xor_cse_481 ^ state_4_4_47_lpi_3
      ^ state_4_4_54_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_24_sva_1;
  assign state_xor_919_nl = (key3[16]) ^ xor_cse_1776 ^ xor_cse_1778 ^ xor_cse_1801;
  assign state_xor_920_nl = xor_cse_57 ^ xor_cse_201 ^ xor_cse_490 ^ state_4_4_48_lpi_3
      ^ state_4_4_55_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_25_sva_1;
  assign state_xor_921_nl = (key3[17]) ^ xor_cse_1773 ^ xor_cse_1781 ^ xor_cse_1799;
  assign state_xor_922_nl = xor_cse_73 ^ xor_cse_214 ^ xor_cse_500 ^ xor_cse_753;
  assign state_xor_923_nl = (key3[18]) ^ xor_cse_1785 ^ xor_cse_1768 ^ xor_cse_1797;
  assign state_xor_924_nl = xor_cse_85 ^ xor_cse_224 ^ xor_cse_516 ^ state_4_4_50_lpi_3
      ^ state_4_4_57_lpi_3 ^ state_1_1_31_0_lpi_4_27;
  assign state_xor_925_nl = (key3[19]) ^ xor_cse_1789 ^ xor_cse_1763 ^ xor_cse_1795;
  assign state_xor_926_nl = xor_cse_100 ^ xor_cse_1 ^ xor_cse_522 ^ xor_cse_763;
  assign state_xor_927_nl = (key3[20]) ^ xor_cse_1792 ^ xor_cse_1758 ^ xor_cse_1793;
  assign state_xor_928_nl = xor_cse_15 ^ xor_cse_526 ^ xor_cse_2903 ^ state_4_4_52_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1 ^ Encrypt_Top_sbox_2_and_2_cse_29_sva_1;
  assign state_xor_929_nl = (key3[21]) ^ xor_cse_1078 ^ xor_cse_1787 ^ xor_cse_1788;
  assign state_xor_930_nl = xor_cse_29 ^ xor_cse_2906 ^ state_4_4_53_lpi_3 ^ state_3_60_lpi_3
      ^ Encrypt_Top_sbox_1_and_cse_30_sva_1 ^ state_4_4_30_lpi_3 ^ xor_cse_775;
  assign state_xor_931_nl = (key3[22]) ^ xor_cse_1087 ^ xor_cse_1783 ^ xor_cse_1784;
  assign state_xor_932_nl = xor_cse_44 ^ xor_cse_536 ^ xor_cse_2909 ^ state_4_4_54_lpi_3
      ^ state_3_61_lpi_3 ^ Encrypt_Top_sbox_2_and_2_cse_31_sva_1;
  assign state_xor_933_nl = (key3[23]) ^ xor_cse_1097 ^ xor_cse_1778 ^ xor_cse_1779;
  assign state_xor_934_nl = xor_cse_57 ^ xor_cse_4 ^ xor_cse_2912 ^ state_4_4_55_lpi_3
      ^ state_1_1_63_32_lpi_4_30 ^ state_4_4_32_lpi_3;
  assign state_xor_935_nl = (key3[24]) ^ xor_cse_1773 ^ xor_cse_1732 ^ xor_cse_1774;
  assign state_xor_936_nl = xor_cse_42 ^ xor_cse_73 ^ xor_cse_18 ^ xor_cse_794;
  assign state_xor_937_nl = (key3[25]) ^ xor_cse_1738 ^ xor_cse_1768 ^ xor_cse_1769;
  assign state_xor_938_nl = xor_cse_56 ^ xor_cse_85 ^ xor_cse_30 ^ xor_cse_801;
  assign state_xor_939_nl = (key3[26]) ^ xor_cse_1745 ^ xor_cse_1763 ^ xor_cse_1764;
  assign state_xor_940_nl = xor_cse_70 ^ xor_cse_100 ^ xor_cse_46 ^ xor_cse_2426;
  assign state_xor_941_nl = (key3[27]) ^ xor_cse_1752 ^ xor_cse_1758 ^ xor_cse_1759;
  assign state_xor_942_nl = xor_cse_84 ^ xor_cse_59 ^ xor_cse_2903 ^ Encrypt_Top_sbox_2_and_2_cse_59_sva_1
      ^ state_4_4_2_lpi_3 ^ state_4_4_36_lpi_3;
  assign state_xor_943_nl = (key3[28]) ^ xor_cse_1078 ^ xor_cse_1753 ^ xor_cse_1754;
  assign state_xor_944_nl = state_3_60_lpi_3 ^ xor_cse_74 ^ xor_cse_2906 ^ xor_cse_2184;
  assign state_xor_945_nl = (key3[29]) ^ xor_cse_1087 ^ xor_cse_1746 ^ xor_cse_1747;
  assign state_xor_946_nl = xor_cse_111 ^ xor_cse_87 ^ xor_cse_2909 ^ state_3_61_lpi_3
      ^ state_4_4_4_lpi_3 ^ state_4_4_38_lpi_3;
  assign state_xor_947_nl = (key3[30]) ^ xor_cse_1739 ^ xor_cse_1097 ^ xor_cse_1740;
  assign state_xor_948_nl = state_1_1_63_32_lpi_4_30 ^ xor_cse_98 ^ xor_cse_2912
      ^ xor_cse_2221;
  assign state_xor_949_nl = (key3[31]) ^ xor_cse_1731 ^ xor_cse_1732 ^ xor_cse_1733;
  assign state_xor_950_nl = xor_cse_136 ^ xor_cse_42 ^ xor_cse_113 ^ xor_cse_2241;
  assign state_xor_951_nl = (key4[8]) ^ xor_cse_1781 ^ xor_cse_1743 ^ xor_cse_1782;
  assign state_xor_952_nl = xor_cse_214 ^ xor_cse_159 ^ xor_cse_673 ^ xor_cse_854;
  assign state_xor_953_nl = (key4[9]) ^ xor_cse_1785 ^ xor_cse_1750 ^ xor_cse_1786;
  assign state_xor_954_nl = xor_cse_170 ^ xor_cse_224 ^ xor_cse_469 ^ state_4_4_9_lpi_3
      ^ Encrypt_Top_sbox_2_and_2_cse_16_sva_1 ^ state_4_4_50_lpi_3;
  assign state_xor_685_nl = (key2[10]) ^ xor_cse_1845 ^ xor_cse_1904 ^ xor_cse_1963;
  assign state_xor_686_nl = (key2[11]) ^ xor_cse_1868 ^ xor_cse_1916 ^ xor_cse_1970;
  assign state_xor_687_nl = (key2[12]) ^ xor_cse_1886 ^ xor_cse_1922 ^ xor_cse_1976;
  assign state_xor_688_nl = (key2[13]) ^ xor_cse_1895 ^ xor_cse_1928 ^ xor_cse_1982;
  assign state_xor_689_nl = (key2[14]) ^ xor_cse_1877 ^ xor_cse_1936 ^ xor_cse_1988;
  assign state_xor_871_nl = xor_cse_1738 ^ xor_cse_379 ^ xor_cse_403 ^ (key4[23])
      ^ state_4_3_31_0_sva_23 ^ state_4_3_31_0_sva_30 ^ Encrypt_Top_sbox_and_2_cse_0_sva_1;
  assign state_xor_872_nl = xor_cse_1745 ^ xor_cse_390 ^ xor_cse_415 ^ (key4[24])
      ^ state_4_3_31_0_sva_24 ^ state_4_3_31_0_sva_31 ^ Encrypt_Top_sbox_and_2_cse_1_sva_1;
  assign state_xnor_176_nl = ~(xor_cse_806 ^ xor_cse_813 ^ xor_cse_1301 ^ state_2_0_1_lpi_6
      ^ state_2_1_1_lpi_6 ^ state_2_6_1_lpi_6);
  assign state_xnor_177_nl = ~(xor_cse_813 ^ xor_cse_821 ^ xor_cse_1311 ^ state_2_1_1_lpi_6
      ^ state_2_2_1_lpi_6 ^ state_2_7_1_lpi_6);
  assign state_xnor_178_nl = ~(xor_cse_821 ^ xor_cse_826 ^ xor_cse_850 ^ state_2_2_1_lpi_6
      ^ state_2_3_1_lpi_6);
  assign state_xnor_179_nl = ~(xor_cse_826 ^ xor_cse_833 ^ xor_cse_851 ^ state_2_3_1_lpi_6
      ^ state_2_4_1_lpi_6);
  assign state_xnor_180_nl = ~(xor_cse_465 ^ xor_cse_833 ^ xor_cse_839 ^ state_2_4_1_lpi_6
      ^ state_2_5_1_lpi_6);
  assign state_xnor_181_nl = ~(xor_cse_839 ^ xor_cse_1301 ^ xor_cse_466 ^ state_2_5_1_lpi_6
      ^ state_2_6_1_lpi_6);
  assign state_xnor_182_nl = ~(xor_cse_1301 ^ xor_cse_1311 ^ xor_cse_477 ^ state_2_6_1_lpi_6
      ^ state_2_7_1_lpi_6);
  assign state_xnor_183_nl = ~(state_2_7_1_lpi_6 ^ xor_cse_1311 ^ xor_cse_850 ^ xor_cse_488);
  assign operator_8_false_mux_1_nl = MUX_v_8_2_2(adlen, plen, fsm_output[13]);
  assign nl_z_out = conv_u2u_8_9(operator_8_false_mux_1_nl) + 9'b111111111;
  assign z_out = nl_z_out[8:0];
  assign AD_P6_mux_2_nl = MUX_v_2_2_2((AD_P6_j_2_0_sva_2[2:1]), (z_out_2[3:2]), or_1265_cse);
  assign nl_AD_P6_acc_nl = ({1'b1 , AD_P6_mux_2_nl}) + 3'b001;
  assign AD_P6_acc_nl = nl_AD_P6_acc_nl[2:0];
  assign z_out_1_2 = readslicef_3_1_2(AD_P6_acc_nl);
  assign or_2257_nl = (fsm_output[13]) | (fsm_output[5]);
  assign INIT_P12_mux_2_nl = MUX_v_3_2_2((signext_3_1(ADLEN_i_7_0_sva_3_0[3])), ADLEN_i_7_0_sva_6_4,
      or_2257_nl);
  assign nl_z_out_2 = conv_u2u_7_8({INIT_P12_mux_2_nl , ADLEN_i_7_0_sva_3_0}) + 8'b00000001;
  assign z_out_2 = nl_z_out_2[7:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_3_1_2;
    input [2:0] vector;
    reg [2:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_3_1_2 = tmp[0:0];
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input  vector;
  begin
    signext_3_1= {{2{vector}}, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_2_3 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_3 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Encrypt_Top
// ------------------------------------------------------------------


module Encrypt_Top (
  clk, rst, arst_n, key1, key2, key3, key4, nonce1, nonce2, nonce3, nonce4, adlen,
      plen, data_in_rsc_dat, data_in_rsc_vld, data_in_rsc_rdy, data_out_rsc_dat,
      data_out_rsc_vld, data_out_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [31:0] key1;
  input [31:0] key2;
  input [31:0] key3;
  input [31:0] key4;
  input [31:0] nonce1;
  input [31:0] nonce2;
  input [31:0] nonce3;
  input [31:0] nonce4;
  input [7:0] adlen;
  input [7:0] plen;
  input [31:0] data_in_rsc_dat;
  input data_in_rsc_vld;
  output data_in_rsc_rdy;
  output [31:0] data_out_rsc_dat;
  output data_out_rsc_vld;
  input data_out_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  Encrypt_Top_run Encrypt_Top_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .key1(key1),
      .key2(key2),
      .key3(key3),
      .key4(key4),
      .nonce1(nonce1),
      .nonce2(nonce2),
      .nonce3(nonce3),
      .nonce4(nonce4),
      .adlen(adlen),
      .plen(plen),
      .data_in_rsc_dat(data_in_rsc_dat),
      .data_in_rsc_vld(data_in_rsc_vld),
      .data_in_rsc_rdy(data_in_rsc_rdy),
      .data_out_rsc_dat(data_out_rsc_dat),
      .data_out_rsc_vld(data_out_rsc_vld),
      .data_out_rsc_rdy(data_out_rsc_rdy)
    );
endmodule



