
//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ../ATTENTION_IP_Attention_Calculator.v4/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   b08092@cad29.ee.ntu.edu.tw
//  Generated date: Wed Jun 12 20:29:13 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, LOOPL1_C_0_tr0, LOOPL1_C_0_tr1, LOOPK2_C_0_tr0,
      LOOPK3_C_0_tr0, LOOPL2_C_0_tr0, LOOPK4_C_1_tr0, LOOPK5_C_1_tr0, LOOPJ1_C_3_tr0,
      LOOPI1_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [16:0] fsm_output;
  reg [16:0] fsm_output;
  input LOOPL1_C_0_tr0;
  input LOOPL1_C_0_tr1;
  input LOOPK2_C_0_tr0;
  input LOOPK3_C_0_tr0;
  input LOOPL2_C_0_tr0;
  input LOOPK4_C_1_tr0;
  input LOOPK5_C_1_tr0;
  input LOOPJ1_C_3_tr0;
  input LOOPI1_C_0_tr0;


  // FSM State Type Declaration for ATTENTION_IP_Attention_Calculator_run_run_fsm_1
  parameter
    main_C_0 = 5'd0,
    LOOPJ1_C_0 = 5'd1,
    LOOPK1_C_0 = 5'd2,
    LOOPL1_C_0 = 5'd3,
    LOOPK1_C_1 = 5'd4,
    LOOPK2_C_0 = 5'd5,
    LOOPJ1_C_1 = 5'd6,
    LOOPK3_C_0 = 5'd7,
    LOOPJ1_C_2 = 5'd8,
    LOOPK4_C_0 = 5'd9,
    LOOPL2_C_0 = 5'd10,
    LOOPK4_C_1 = 5'd11,
    LOOPK5_C_0 = 5'd12,
    LOOPK5_C_1 = 5'd13,
    LOOPJ1_C_3 = 5'd14,
    LOOPI1_C_0 = 5'd15,
    main_C_1 = 5'd16;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ATTENTION_IP_Attention_Calculator_run_run_fsm_1
    case (state_var)
      LOOPJ1_C_0 : begin
        fsm_output = 17'b00000000000000010;
        state_var_NS = LOOPK1_C_0;
      end
      LOOPK1_C_0 : begin
        fsm_output = 17'b00000000000000100;
        state_var_NS = LOOPL1_C_0;
      end
      LOOPL1_C_0 : begin
        fsm_output = 17'b00000000000001000;
        if ( LOOPL1_C_0_tr0 ) begin
          state_var_NS = LOOPK2_C_0;
        end
        else if ( LOOPL1_C_0_tr1 ) begin
          state_var_NS = LOOPL1_C_0;
        end
        else begin
          state_var_NS = LOOPK1_C_1;
        end
      end
      LOOPK1_C_1 : begin
        fsm_output = 17'b00000000000010000;
        state_var_NS = LOOPK1_C_0;
      end
      LOOPK2_C_0 : begin
        fsm_output = 17'b00000000000100000;
        if ( LOOPK2_C_0_tr0 ) begin
          state_var_NS = LOOPJ1_C_1;
        end
        else begin
          state_var_NS = LOOPK2_C_0;
        end
      end
      LOOPJ1_C_1 : begin
        fsm_output = 17'b00000000001000000;
        state_var_NS = LOOPK3_C_0;
      end
      LOOPK3_C_0 : begin
        fsm_output = 17'b00000000010000000;
        if ( LOOPK3_C_0_tr0 ) begin
          state_var_NS = LOOPJ1_C_2;
        end
        else begin
          state_var_NS = LOOPK3_C_0;
        end
      end
      LOOPJ1_C_2 : begin
        fsm_output = 17'b00000000100000000;
        state_var_NS = LOOPK4_C_0;
      end
      LOOPK4_C_0 : begin
        fsm_output = 17'b00000001000000000;
        state_var_NS = LOOPL2_C_0;
      end
      LOOPL2_C_0 : begin
        fsm_output = 17'b00000010000000000;
        if ( LOOPL2_C_0_tr0 ) begin
          state_var_NS = LOOPK4_C_1;
        end
        else begin
          state_var_NS = LOOPL2_C_0;
        end
      end
      LOOPK4_C_1 : begin
        fsm_output = 17'b00000100000000000;
        if ( LOOPK4_C_1_tr0 ) begin
          state_var_NS = LOOPK5_C_0;
        end
        else begin
          state_var_NS = LOOPK4_C_0;
        end
      end
      LOOPK5_C_0 : begin
        fsm_output = 17'b00001000000000000;
        state_var_NS = LOOPK5_C_1;
      end
      LOOPK5_C_1 : begin
        fsm_output = 17'b00010000000000000;
        if ( LOOPK5_C_1_tr0 ) begin
          state_var_NS = LOOPJ1_C_3;
        end
        else begin
          state_var_NS = LOOPK5_C_0;
        end
      end
      LOOPJ1_C_3 : begin
        fsm_output = 17'b00100000000000000;
        if ( LOOPJ1_C_3_tr0 ) begin
          state_var_NS = LOOPI1_C_0;
        end
        else begin
          state_var_NS = LOOPJ1_C_0;
        end
      end
      LOOPI1_C_0 : begin
        fsm_output = 17'b01000000000000000;
        if ( LOOPI1_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = LOOPJ1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 17'b10000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 17'b00000000000000001;
        state_var_NS = LOOPJ1_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_staller
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_staller (
  run_wen, q_chan2_rsci_wen_comp, k_chan2_rsci_wen_comp, v_chan2_rsci_wen_comp, dout_chan_rsci_wen_comp
);
  output run_wen;
  input q_chan2_rsci_wen_comp;
  input k_chan2_rsci_wen_comp;
  input v_chan2_rsci_wen_comp;
  input dout_chan_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = q_chan2_rsci_wen_comp & k_chan2_rsci_wen_comp & v_chan2_rsci_wen_comp
      & dout_chan_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci_dout_chan_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci_dout_chan_wait_ctrl (
  dout_chan_rsci_iswt0, dout_chan_rsci_biwt, dout_chan_rsci_irdy
);
  input dout_chan_rsci_iswt0;
  output dout_chan_rsci_biwt;
  input dout_chan_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign dout_chan_rsci_biwt = dout_chan_rsci_iswt0 & dout_chan_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci_v_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci_v_chan2_wait_ctrl (
  v_chan2_rsci_iswt0, v_chan2_rsci_biwt, v_chan2_rsci_ivld
);
  input v_chan2_rsci_iswt0;
  output v_chan2_rsci_biwt;
  input v_chan2_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign v_chan2_rsci_biwt = v_chan2_rsci_iswt0 & v_chan2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci_k_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci_k_chan2_wait_ctrl (
  k_chan2_rsci_iswt0, k_chan2_rsci_biwt, k_chan2_rsci_ivld
);
  input k_chan2_rsci_iswt0;
  output k_chan2_rsci_biwt;
  input k_chan2_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign k_chan2_rsci_biwt = k_chan2_rsci_iswt0 & k_chan2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci_q_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci_q_chan2_wait_ctrl (
  q_chan2_rsci_iswt0, q_chan2_rsci_biwt, q_chan2_rsci_ivld
);
  input q_chan2_rsci_iswt0;
  output q_chan2_rsci_biwt;
  input q_chan2_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign q_chan2_rsci_biwt = q_chan2_rsci_iswt0 & q_chan2_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci (
  dout_chan_rsc_dat, dout_chan_rsc_vld, dout_chan_rsc_rdy, dout_chan_rsci_oswt, dout_chan_rsci_wen_comp,
      dout_chan_rsci_idat
);
  output [15:0] dout_chan_rsc_dat;
  output dout_chan_rsc_vld;
  input dout_chan_rsc_rdy;
  input dout_chan_rsci_oswt;
  output dout_chan_rsci_wen_comp;
  input [15:0] dout_chan_rsci_idat;


  // Interconnect Declarations
  wire dout_chan_rsci_biwt;
  wire dout_chan_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd7),
  .width(32'sd16)) dout_chan_rsci (
      .irdy(dout_chan_rsci_irdy),
      .ivld(dout_chan_rsci_oswt),
      .idat(dout_chan_rsci_idat),
      .rdy(dout_chan_rsc_rdy),
      .vld(dout_chan_rsc_vld),
      .dat(dout_chan_rsc_dat)
    );
  ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci_dout_chan_wait_ctrl ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci_dout_chan_wait_ctrl_inst
      (
      .dout_chan_rsci_iswt0(dout_chan_rsci_oswt),
      .dout_chan_rsci_biwt(dout_chan_rsci_biwt),
      .dout_chan_rsci_irdy(dout_chan_rsci_irdy)
    );
  assign dout_chan_rsci_wen_comp = (~ dout_chan_rsci_oswt) | dout_chan_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci (
  v_chan2_rsc_dat, v_chan2_rsc_vld, v_chan2_rsc_rdy, v_chan2_rsci_oswt, v_chan2_rsci_wen_comp,
      v_chan2_rsci_idat_mxwt
);
  input [1023:0] v_chan2_rsc_dat;
  input v_chan2_rsc_vld;
  output v_chan2_rsc_rdy;
  input v_chan2_rsci_oswt;
  output v_chan2_rsci_wen_comp;
  output [1023:0] v_chan2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire v_chan2_rsci_biwt;
  wire v_chan2_rsci_ivld;
  wire [1023:0] v_chan2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd1024)) v_chan2_rsci (
      .rdy(v_chan2_rsc_rdy),
      .vld(v_chan2_rsc_vld),
      .dat(v_chan2_rsc_dat),
      .irdy(v_chan2_rsci_oswt),
      .ivld(v_chan2_rsci_ivld),
      .idat(v_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci_v_chan2_wait_ctrl ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci_v_chan2_wait_ctrl_inst
      (
      .v_chan2_rsci_iswt0(v_chan2_rsci_oswt),
      .v_chan2_rsci_biwt(v_chan2_rsci_biwt),
      .v_chan2_rsci_ivld(v_chan2_rsci_ivld)
    );
  assign v_chan2_rsci_idat_mxwt = v_chan2_rsci_idat;
  assign v_chan2_rsci_wen_comp = (~ v_chan2_rsci_oswt) | v_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci (
  k_chan2_rsc_dat, k_chan2_rsc_vld, k_chan2_rsc_rdy, k_chan2_rsci_oswt, k_chan2_rsci_wen_comp,
      k_chan2_rsci_idat_mxwt
);
  input [1023:0] k_chan2_rsc_dat;
  input k_chan2_rsc_vld;
  output k_chan2_rsc_rdy;
  input k_chan2_rsci_oswt;
  output k_chan2_rsci_wen_comp;
  output [1023:0] k_chan2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire k_chan2_rsci_biwt;
  wire k_chan2_rsci_ivld;
  wire [1023:0] k_chan2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd1024)) k_chan2_rsci (
      .rdy(k_chan2_rsc_rdy),
      .vld(k_chan2_rsc_vld),
      .dat(k_chan2_rsc_dat),
      .irdy(k_chan2_rsci_oswt),
      .ivld(k_chan2_rsci_ivld),
      .idat(k_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci_k_chan2_wait_ctrl ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci_k_chan2_wait_ctrl_inst
      (
      .k_chan2_rsci_iswt0(k_chan2_rsci_oswt),
      .k_chan2_rsci_biwt(k_chan2_rsci_biwt),
      .k_chan2_rsci_ivld(k_chan2_rsci_ivld)
    );
  assign k_chan2_rsci_idat_mxwt = k_chan2_rsci_idat;
  assign k_chan2_rsci_wen_comp = (~ k_chan2_rsci_oswt) | k_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci (
  q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy, q_chan2_rsci_oswt, q_chan2_rsci_wen_comp,
      q_chan2_rsci_idat_mxwt
);
  input [1023:0] q_chan2_rsc_dat;
  input q_chan2_rsc_vld;
  output q_chan2_rsc_rdy;
  input q_chan2_rsci_oswt;
  output q_chan2_rsci_wen_comp;
  output [1023:0] q_chan2_rsci_idat_mxwt;


  // Interconnect Declarations
  wire q_chan2_rsci_biwt;
  wire q_chan2_rsci_ivld;
  wire [1023:0] q_chan2_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd4),
  .width(32'sd1024)) q_chan2_rsci (
      .rdy(q_chan2_rsc_rdy),
      .vld(q_chan2_rsc_vld),
      .dat(q_chan2_rsc_dat),
      .irdy(q_chan2_rsci_oswt),
      .ivld(q_chan2_rsci_ivld),
      .idat(q_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci_q_chan2_wait_ctrl ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci_q_chan2_wait_ctrl_inst
      (
      .q_chan2_rsci_iswt0(q_chan2_rsci_oswt),
      .q_chan2_rsci_biwt(q_chan2_rsci_biwt),
      .q_chan2_rsci_ivld(q_chan2_rsci_ivld)
    );
  assign q_chan2_rsci_idat_mxwt = q_chan2_rsci_idat;
  assign q_chan2_rsci_wen_comp = (~ q_chan2_rsci_oswt) | q_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator_run
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator_run (
  clk, rst, arst_n, head, length, dim, q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy,
      k_chan2_rsc_dat, k_chan2_rsc_vld, k_chan2_rsc_rdy, v_chan2_rsc_dat, v_chan2_rsc_vld,
      v_chan2_rsc_rdy, dout_chan_rsc_dat, dout_chan_rsc_vld, dout_chan_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [1023:0] q_chan2_rsc_dat;
  input q_chan2_rsc_vld;
  output q_chan2_rsc_rdy;
  input [1023:0] k_chan2_rsc_dat;
  input k_chan2_rsc_vld;
  output k_chan2_rsc_rdy;
  input [1023:0] v_chan2_rsc_dat;
  input v_chan2_rsc_vld;
  output v_chan2_rsc_rdy;
  output [15:0] dout_chan_rsc_dat;
  output dout_chan_rsc_vld;
  input dout_chan_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire q_chan2_rsci_wen_comp;
  wire [1023:0] q_chan2_rsci_idat_mxwt;
  wire k_chan2_rsci_wen_comp;
  wire [1023:0] k_chan2_rsci_idat_mxwt;
  wire v_chan2_rsci_wen_comp;
  wire [1023:0] v_chan2_rsci_idat_mxwt;
  wire dout_chan_rsci_wen_comp;
  reg [15:0] dout_chan_rsci_idat;
  wire [16:0] fsm_output;
  wire LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp;
  wire LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp;
  wire LOOPK4_LOOPK4_if_1_and_tmp;
  wire LOOPK3_if_unequal_tmp;
  wire LOOPK3_if_equal_tmp;
  wire LOOPL1_LOOPL1_nor_tmp;
  wire LOOPL1_LOOPL1_and_tmp;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire or_dcpl_215;
  wire or_dcpl_216;
  wire or_dcpl_217;
  wire or_dcpl_218;
  wire or_dcpl_219;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire or_dcpl_222;
  wire or_dcpl_223;
  wire or_dcpl_224;
  wire or_dcpl_225;
  wire or_dcpl_226;
  wire and_dcpl_97;
  wire or_dcpl_229;
  wire or_dcpl_230;
  wire and_dcpl_101;
  wire or_dcpl_233;
  wire or_dcpl_234;
  wire or_dcpl_237;
  wire or_dcpl_240;
  wire or_dcpl_243;
  wire or_dcpl_246;
  wire or_dcpl_247;
  wire or_dcpl_248;
  wire and_dcpl_115;
  wire and_dcpl_116;
  wire and_dcpl_118;
  wire and_dcpl_119;
  wire or_dcpl_250;
  wire or_dcpl_251;
  wire or_dcpl_252;
  wire or_dcpl_253;
  wire or_dcpl_254;
  wire and_dcpl_121;
  wire and_dcpl_122;
  wire and_dcpl_124;
  wire and_dcpl_125;
  wire and_dcpl_126;
  wire and_dcpl_127;
  wire or_dcpl_256;
  wire or_dcpl_257;
  wire or_dcpl_258;
  wire or_dcpl_259;
  wire or_dcpl_260;
  wire or_dcpl_261;
  wire and_dcpl_129;
  wire or_dcpl_263;
  wire or_dcpl_264;
  wire and_dcpl_132;
  wire and_dcpl_134;
  wire and_dcpl_135;
  wire or_dcpl_266;
  wire or_dcpl_267;
  wire or_dcpl_268;
  wire or_dcpl_269;
  wire and_dcpl_137;
  wire and_dcpl_139;
  wire or_dcpl_271;
  wire or_dcpl_272;
  wire or_dcpl_273;
  wire and_dcpl_141;
  wire and_dcpl_143;
  wire or_dcpl_275;
  wire or_dcpl_276;
  wire or_dcpl_277;
  wire and_dcpl_145;
  wire or_dcpl_279;
  wire or_dcpl_280;
  wire and_dcpl_148;
  wire or_dcpl_282;
  wire or_dcpl_284;
  wire and_dcpl_154;
  wire or_dcpl_286;
  wire or_dcpl_287;
  wire or_dcpl_289;
  wire and_dcpl_159;
  wire or_dcpl_291;
  wire or_dcpl_292;
  wire or_dcpl_294;
  wire or_dcpl_296;
  wire or_dcpl_298;
  wire or_dcpl_300;
  wire or_dcpl_301;
  wire and_dcpl_169;
  wire and_dcpl_171;
  wire or_dcpl_303;
  wire or_dcpl_304;
  wire or_dcpl_305;
  wire and_dcpl_173;
  wire and_dcpl_175;
  wire or_dcpl_307;
  wire or_dcpl_308;
  wire or_dcpl_309;
  wire and_dcpl_177;
  wire or_dcpl_311;
  wire or_dcpl_312;
  wire and_dcpl_180;
  wire or_dcpl_314;
  wire or_dcpl_315;
  wire and_dcpl_183;
  wire or_dcpl_317;
  wire or_dcpl_318;
  wire and_dcpl_186;
  wire or_dcpl_320;
  wire or_dcpl_321;
  wire and_dcpl_189;
  wire or_dcpl_323;
  wire or_dcpl_324;
  wire and_dcpl_192;
  wire or_dcpl_326;
  wire or_dcpl_328;
  wire or_dcpl_330;
  wire or_dcpl_332;
  wire or_dcpl_334;
  wire or_dcpl_336;
  wire or_dcpl_338;
  wire or_dcpl_340;
  wire or_dcpl_342;
  wire or_dcpl_343;
  wire and_dcpl_211;
  wire or_dcpl_345;
  wire or_dcpl_346;
  wire and_dcpl_214;
  wire or_dcpl_348;
  wire or_dcpl_350;
  wire or_dcpl_352;
  wire or_dcpl_354;
  wire or_dcpl_356;
  wire or_dcpl_358;
  wire or_dcpl_360;
  wire or_dcpl_362;
  wire or_dcpl_364;
  wire or_dcpl_366;
  wire or_dcpl_368;
  wire or_dcpl_370;
  wire or_dcpl_372;
  wire or_dcpl_374;
  wire or_dcpl_376;
  wire and_dcpl_245;
  wire and_dcpl_246;
  wire and_dcpl_247;
  wire and_dcpl_248;
  wire and_dcpl_251;
  wire and_dcpl_252;
  wire and_dcpl_253;
  wire and_dcpl_254;
  wire and_dcpl_256;
  wire and_dcpl_258;
  wire and_dcpl_264;
  wire and_dcpl_265;
  wire and_dcpl_267;
  wire and_dcpl_268;
  wire and_dcpl_276;
  wire and_dcpl_278;
  wire and_dcpl_286;
  wire and_dcpl_288;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_300;
  wire and_dcpl_301;
  wire and_dcpl_303;
  wire and_dcpl_305;
  wire and_dcpl_348;
  wire or_tmp_553;
  wire and_363_cse;
  wire and_671_cse;
  reg LOOPK1_endflag_sva;
  reg [31:0] LOOPL2_l_sva;
  wire LOOPK3_and_stg_3_15_sva_1;
  wire LOOPK3_and_stg_3_1_sva_1;
  wire LOOPK3_and_stg_3_14_sva_1;
  wire LOOPK3_and_stg_3_2_sva_1;
  wire LOOPK3_and_stg_3_13_sva_1;
  wire LOOPK3_and_stg_3_3_sva_1;
  wire LOOPK3_and_stg_3_12_sva_1;
  wire LOOPK3_and_stg_3_4_sva_1;
  wire LOOPK3_and_stg_3_11_sva_1;
  wire LOOPK3_and_stg_3_5_sva_1;
  wire LOOPK3_and_stg_3_10_sva_1;
  wire LOOPK3_and_stg_3_6_sva_1;
  wire LOOPK3_and_stg_3_9_sva_1;
  wire LOOPK3_and_stg_3_7_sva_1;
  wire LOOPK3_and_stg_3_8_sva_1;
  wire LOOPK3_and_stg_2_0_sva_1;
  wire LOOPK3_and_stg_2_1_sva_1;
  wire LOOPK3_and_stg_2_2_sva_1;
  wire LOOPK3_and_stg_2_3_sva_1;
  wire LOOPK3_and_stg_2_4_sva_1;
  wire LOOPK3_and_stg_2_5_sva_1;
  wire LOOPK3_and_stg_2_6_sva_1;
  wire LOOPK3_and_stg_2_7_sva_1;
  wire LOOPK3_and_stg_1_0_sva_1;
  wire LOOPK3_and_stg_1_1_sva_1;
  wire LOOPK3_and_stg_1_2_sva_1;
  wire LOOPK3_and_stg_1_3_sva_1;
  wire LOOPK2_and_115_cse_sva_1;
  wire LOOPK2_else_or_tmp_3;
  wire LOOPK2_else_or_tmp_2;
  wire LOOPK2_and_113_cse_sva_1;
  wire LOOPK2_and_111_cse_sva_1;
  wire LOOPK2_and_109_cse_sva_1;
  wire LOOPK2_and_107_cse_sva_1;
  wire LOOPK2_and_105_cse_sva_1;
  wire LOOPK2_and_103_cse_sva_1;
  wire LOOPK2_and_101_cse_sva_1;
  wire LOOPK2_and_99_cse_sva_1;
  wire LOOPK2_and_97_cse_sva_1;
  wire LOOPK2_and_95_cse_sva_1;
  wire LOOPK2_and_93_cse_sva_1;
  wire LOOPK2_and_91_cse_sva_1;
  wire LOOPK2_and_89_cse_sva_1;
  wire LOOPK2_and_87_cse_sva_1;
  wire LOOPK2_and_85_cse_sva_1;
  wire LOOPK2_and_83_cse_sva_1;
  wire LOOPK2_and_81_cse_sva_1;
  wire LOOPK2_and_79_cse_sva_1;
  wire LOOPK2_and_77_cse_sva_1;
  wire LOOPK2_and_75_cse_sva_1;
  wire LOOPK2_and_73_cse_sva_1;
  wire LOOPK2_and_71_cse_sva_1;
  wire LOOPK2_and_69_cse_sva_1;
  wire LOOPK2_and_67_cse_sva_1;
  wire LOOPK2_and_65_cse_sva_1;
  wire LOOPK2_and_63_cse_sva_1;
  wire LOOPK2_and_61_cse_sva_1;
  wire LOOPK2_and_60_cse_sva_1;
  wire LOOPK2_and_62_cse_sva_1;
  wire LOOPK2_and_64_cse_sva_1;
  wire LOOPK2_and_66_cse_sva_1;
  wire LOOPK2_and_68_cse_sva_1;
  wire LOOPK2_and_70_cse_sva_1;
  wire LOOPK2_and_72_cse_sva_1;
  wire LOOPK2_and_74_cse_sva_1;
  wire LOOPK2_and_76_cse_sva_1;
  wire LOOPK2_and_78_cse_sva_1;
  wire LOOPK2_and_80_cse_sva_1;
  wire LOOPK2_and_82_cse_sva_1;
  wire LOOPK2_and_84_cse_sva_1;
  wire LOOPK2_and_86_cse_sva_1;
  wire LOOPK2_and_88_cse_sva_1;
  wire LOOPK2_and_90_cse_sva_1;
  wire LOOPK2_and_92_cse_sva_1;
  wire LOOPK2_and_94_cse_sva_1;
  wire LOOPK2_and_96_cse_sva_1;
  wire LOOPK2_and_98_cse_sva_1;
  wire LOOPK2_and_100_cse_sva_1;
  wire LOOPK2_and_102_cse_sva_1;
  wire LOOPK2_and_104_cse_sva_1;
  wire LOOPK2_and_106_cse_sva_1;
  wire LOOPK2_and_108_cse_sva_1;
  wire LOOPK2_and_110_cse_sva_1;
  wire LOOPK2_and_112_cse_sva_1;
  wire LOOPK2_and_114_cse_sva_1;
  wire LOOPK2_and_stg_4_23_sva_1;
  wire LOOPK2_and_stg_4_0_sva_1;
  wire LOOPK2_and_stg_4_22_sva_1;
  wire LOOPK2_and_stg_4_1_sva_1;
  wire LOOPK2_and_stg_4_21_sva_1;
  wire LOOPK2_and_stg_4_2_sva_1;
  wire LOOPK2_and_stg_4_20_sva_1;
  wire LOOPK2_and_stg_4_3_sva_1;
  wire LOOPK2_and_stg_4_19_sva_1;
  wire LOOPK2_and_stg_4_4_sva_1;
  wire LOOPK2_and_stg_4_18_sva_1;
  wire LOOPK2_and_stg_4_5_sva_1;
  wire LOOPK2_and_stg_4_17_sva_1;
  wire LOOPK2_and_stg_4_6_sva_1;
  wire LOOPK2_and_stg_4_16_sva_1;
  wire LOOPK2_and_stg_4_7_sva_1;
  wire LOOPK2_and_stg_4_15_sva_1;
  wire LOOPK2_and_stg_4_8_sva_1;
  wire LOOPK2_and_stg_4_14_sva_1;
  wire LOOPK2_and_stg_4_9_sva_1;
  wire LOOPK2_and_stg_4_13_sva_1;
  wire LOOPK2_and_stg_4_10_sva_1;
  wire LOOPK2_and_stg_4_12_sva_1;
  wire LOOPK2_and_stg_4_11_sva_1;
  wire LOOPK2_and_stg_3_0_sva_1;
  wire LOOPK1_and_stg_3_11_sva_1;
  wire LOOPK1_and_stg_2_0_sva_1;
  wire LOOPK1_and_stg_2_1_sva_1;
  wire LOOPK1_and_stg_2_2_sva_1;
  wire LOOPK1_and_stg_2_3_sva_1;
  wire LOOPK1_and_stg_2_4_sva_1;
  wire LOOPK1_and_stg_2_5_sva_1;
  wire LOOPK1_and_stg_2_6_sva_1;
  wire LOOPK1_and_stg_2_7_sva_1;
  wire LOOPK1_and_stg_1_0_sva_1;
  wire LOOPK1_and_stg_1_1_sva_1;
  wire LOOPK1_and_stg_1_2_sva_1;
  wire LOOPK1_and_stg_1_3_sva_1;
  reg [7:0] cnt_sva;
  reg LOOPK1_and_60_itm;
  reg LOOPK1_slc_cnt_5_0_10_itm;
  reg LOOPK1_and_stg_3_12_sva;
  reg LOOPK1_slc_cnt_5_0_66_itm;
  reg LOOPK1_and_stg_3_10_sva;
  reg LOOPK1_and_stg_3_13_sva;
  reg LOOPK1_and_stg_3_9_sva;
  reg LOOPK1_and_stg_3_14_sva;
  reg LOOPK1_and_stg_3_8_sva;
  reg LOOPK1_and_stg_3_15_sva;
  reg LOOPK1_and_stg_2_7_sva;
  reg LOOPK1_slc_cnt_5_0_9_itm;
  reg LOOPK1_and_stg_2_0_sva;
  reg LOOPK1_and_stg_2_6_sva;
  reg LOOPK1_and_stg_2_1_sva;
  reg LOOPK1_and_stg_2_5_sva;
  reg LOOPK1_and_stg_2_2_sva;
  reg LOOPK1_and_stg_2_4_sva;
  reg LOOPK1_and_stg_2_3_sva;
  reg LOOPK1_and_stg_3_11_sva;
  wire [37:0] sum_array_0_sva_2_mx0;
  wire [37:0] sum_array_1_sva_2_mx0;
  wire [37:0] sum_array_2_sva_2_mx0;
  wire [37:0] sum_array_3_sva_2_mx0;
  wire [37:0] sum_array_4_sva_2_mx0;
  wire [37:0] sum_array_5_sva_2_mx0;
  wire [37:0] sum_array_6_sva_2_mx0;
  wire [37:0] sum_array_7_sva_2_mx0;
  wire [37:0] sum_array_8_sva_2_mx0;
  wire [37:0] sum_array_9_sva_2_mx0;
  wire [37:0] sum_array_10_sva_2_mx0;
  wire [37:0] sum_array_11_sva_2_mx0;
  wire [37:0] sum_array_12_sva_2_mx0;
  wire [37:0] sum_array_13_sva_2_mx0;
  wire [37:0] sum_array_14_sva_2_mx0;
  wire [37:0] sum_array_15_sva_2_mx0;
  wire [37:0] sum_array_16_sva_2_mx0;
  wire [37:0] sum_array_17_sva_2_mx0;
  wire [37:0] sum_array_18_sva_2_mx0;
  wire [37:0] sum_array_19_sva_2_mx0;
  wire [37:0] sum_array_20_sva_2_mx0;
  wire [37:0] sum_array_21_sva_2_mx0;
  wire [37:0] sum_array_22_sva_2_mx0;
  wire [37:0] sum_array_23_sva_2_mx0;
  wire [37:0] sum_array_24_sva_2_mx0;
  wire [37:0] sum_array_25_sva_2_mx0;
  wire [37:0] sum_array_26_sva_2_mx0;
  wire [37:0] sum_array_27_sva_2_mx0;
  wire [37:0] sum_array_28_sva_2_mx0;
  wire [37:0] sum_array_29_sva_2_mx0;
  wire [37:0] sum_array_30_sva_2_mx0;
  wire [37:0] sum_array_31_sva_2_mx0;
  wire [37:0] sum_array_32_sva_2_mx0;
  wire [37:0] sum_array_33_sva_2_mx0;
  wire [37:0] sum_array_34_sva_2_mx0;
  wire [37:0] sum_array_35_sva_2_mx0;
  wire [37:0] sum_array_36_sva_2_mx0;
  wire [37:0] sum_array_37_sva_2_mx0;
  wire [37:0] sum_array_38_sva_2_mx0;
  wire [37:0] sum_array_39_sva_2_mx0;
  wire [37:0] sum_array_40_sva_2_mx0;
  wire [37:0] sum_array_41_sva_2_mx0;
  wire [37:0] sum_array_42_sva_2_mx0;
  wire [37:0] sum_array_43_sva_2_mx0;
  wire [37:0] sum_array_44_sva_2_mx0;
  wire [37:0] sum_array_45_sva_2_mx0;
  wire [37:0] sum_array_46_sva_2_mx0;
  wire [37:0] sum_array_47_sva_2_mx0;
  wire [37:0] sum_array_48_sva_2_mx0;
  wire [37:0] sum_array_49_sva_2_mx0;
  wire [37:0] sum_array_50_sva_2_mx0;
  wire [37:0] sum_array_51_sva_2_mx0;
  wire [37:0] sum_array_52_sva_2_mx0;
  wire [37:0] sum_array_53_sva_2_mx0;
  wire [37:0] sum_array_54_sva_2_mx0;
  wire [37:0] sum_array_55_sva_2_mx0;
  wire LOOPK2_else_equal_tmp_16;
  wire LOOPK2_else_equal_tmp_130;
  wire LOOPK2_else_equal_tmp_244;
  wire LOOPK2_else_equal_tmp_358;
  wire LOOPK2_else_equal_tmp_472;
  wire LOOPK2_else_equal_tmp_586;
  wire LOOPK2_else_equal_tmp_700;
  wire LOOPK2_else_equal_tmp_814;
  wire LOOPK2_else_equal_tmp_928;
  wire LOOPK2_else_equal_tmp_1042;
  wire LOOPK2_else_equal_tmp_1156;
  wire LOOPK2_else_equal_tmp_1270;
  wire LOOPK2_else_equal_tmp_1384;
  wire LOOPK2_else_equal_tmp_1498;
  wire LOOPK2_else_equal_tmp_1612;
  wire LOOPK2_else_equal_tmp_1726;
  reg reg_q_chan2_rsci_oswt_cse;
  reg reg_k_chan2_rsci_oswt_cse;
  reg reg_v_chan2_rsci_oswt_cse;
  reg reg_dout_chan_rsci_oswt_cse;
  wire LOOPK5_k_nor_seb;
  reg LOOPK5_k_sva_6;
  reg [5:0] LOOPK5_k_sva_5_0;
  wire LOOPL1_if_1_unequal_1_itm;
  wire [5:0] z_out;
  wire [6:0] nl_z_out;
  wire [8:0] z_out_1;
  wire [9:0] nl_z_out_1;
  wire [7:0] z_out_2;
  wire [8:0] nl_z_out_2;
  wire [15:0] z_out_3;
  wire [16:0] nl_z_out_3;
  wire [15:0] z_out_4;
  wire [15:0] z_out_5;
  wire [37:0] z_out_6;
  wire signed [55:0] nl_z_out_6;
  reg [3:0] LOOPI1_i_sva;
  reg [37:0] sum_array_27_lpi_3;
  reg [37:0] sum_array_28_lpi_3;
  reg [37:0] sum_array_26_lpi_3;
  reg [37:0] sum_array_29_lpi_3;
  reg [37:0] sum_array_25_lpi_3;
  reg [37:0] sum_array_30_lpi_3;
  reg [37:0] sum_array_24_lpi_3;
  reg [37:0] sum_array_31_lpi_3;
  reg [37:0] sum_array_23_lpi_3;
  reg [37:0] sum_array_32_lpi_3;
  reg [37:0] sum_array_22_lpi_3;
  reg [37:0] sum_array_33_lpi_3;
  reg [37:0] sum_array_21_lpi_3;
  reg [37:0] sum_array_34_lpi_3;
  reg [37:0] sum_array_20_lpi_3;
  reg [37:0] sum_array_35_lpi_3;
  reg [37:0] sum_array_19_lpi_3;
  reg [37:0] sum_array_36_lpi_3;
  reg [37:0] sum_array_18_lpi_3;
  reg [37:0] sum_array_37_lpi_3;
  reg [37:0] sum_array_17_lpi_3;
  reg [37:0] sum_array_38_lpi_3;
  reg [37:0] sum_array_16_lpi_3;
  reg [37:0] sum_array_39_lpi_3;
  reg [37:0] sum_array_15_lpi_3;
  reg [37:0] sum_array_40_lpi_3;
  reg [37:0] sum_array_14_lpi_3;
  reg [37:0] sum_array_41_lpi_3;
  reg [37:0] sum_array_13_lpi_3;
  reg [37:0] sum_array_42_lpi_3;
  reg [37:0] sum_array_12_lpi_3;
  reg [37:0] sum_array_43_lpi_3;
  reg [37:0] sum_array_11_lpi_3;
  reg [37:0] sum_array_44_lpi_3;
  reg [37:0] sum_array_10_lpi_3;
  reg [37:0] sum_array_45_lpi_3;
  reg [37:0] sum_array_9_lpi_3;
  reg [37:0] sum_array_46_lpi_3;
  reg [37:0] sum_array_8_lpi_3;
  reg [37:0] sum_array_47_lpi_3;
  reg [37:0] sum_array_7_lpi_3;
  reg [37:0] sum_array_48_lpi_3;
  reg [37:0] sum_array_6_lpi_3;
  reg [37:0] sum_array_49_lpi_3;
  reg [37:0] sum_array_5_lpi_3;
  reg [37:0] sum_array_50_lpi_3;
  reg [37:0] sum_array_4_lpi_3;
  reg [37:0] sum_array_51_lpi_3;
  reg [37:0] sum_array_3_lpi_3;
  reg [37:0] sum_array_52_lpi_3;
  reg [37:0] sum_array_2_lpi_3;
  reg [37:0] sum_array_53_lpi_3;
  reg [37:0] sum_array_1_lpi_3;
  reg [37:0] sum_array_54_lpi_3;
  reg [37:0] sum_array_0_lpi_3;
  reg [37:0] sum_array_55_lpi_3;
  reg [15:0] data_out_32_lpi_3;
  reg [15:0] data_out_30_lpi_3;
  reg [15:0] data_out_34_lpi_3;
  reg [15:0] data_out_28_lpi_3;
  reg [15:0] data_out_36_lpi_3;
  reg [15:0] data_out_26_lpi_3;
  reg [15:0] data_out_38_lpi_3;
  reg [15:0] data_out_24_lpi_3;
  reg [15:0] data_out_40_lpi_3;
  reg [15:0] data_out_22_lpi_3;
  reg [15:0] data_out_42_lpi_3;
  reg [15:0] data_out_20_lpi_3;
  reg [15:0] data_out_44_lpi_3;
  reg [15:0] data_out_18_lpi_3;
  reg [15:0] data_out_46_lpi_3;
  reg [15:0] data_out_16_lpi_3;
  reg [15:0] data_out_48_lpi_3;
  reg [15:0] data_out_14_lpi_3;
  reg [15:0] data_out_50_lpi_3;
  reg [15:0] data_out_12_lpi_3;
  reg [15:0] data_out_52_lpi_3;
  reg [15:0] data_out_10_lpi_3;
  reg [15:0] data_out_54_lpi_3;
  reg [15:0] data_out_8_lpi_3;
  reg [15:0] data_out_56_lpi_3;
  reg [15:0] data_out_6_lpi_3;
  reg [15:0] data_out_58_lpi_3;
  reg [15:0] data_out_4_lpi_3;
  reg [15:0] data_out_60_lpi_3;
  reg [15:0] data_out_2_lpi_3;
  reg [15:0] data_out_62_lpi_3;
  reg [15:0] data_out_31_lpi_3;
  reg [15:0] data_out_33_lpi_3;
  reg [15:0] data_out_29_lpi_3;
  reg [15:0] data_out_35_lpi_3;
  reg [15:0] data_out_27_lpi_3;
  reg [15:0] data_out_37_lpi_3;
  reg [15:0] data_out_25_lpi_3;
  reg [15:0] data_out_39_lpi_3;
  reg [15:0] data_out_23_lpi_3;
  reg [15:0] data_out_41_lpi_3;
  reg [15:0] data_out_21_lpi_3;
  reg [15:0] data_out_43_lpi_3;
  reg [15:0] data_out_19_lpi_3;
  reg [15:0] data_out_45_lpi_3;
  reg [15:0] data_out_17_lpi_3;
  reg [15:0] data_out_47_lpi_3;
  reg [15:0] data_out_15_lpi_3;
  reg [15:0] data_out_49_lpi_3;
  reg [15:0] data_out_13_lpi_3;
  reg [15:0] data_out_51_lpi_3;
  reg [15:0] data_out_11_lpi_3;
  reg [15:0] data_out_53_lpi_3;
  reg [15:0] data_out_9_lpi_3;
  reg [15:0] data_out_55_lpi_3;
  reg [15:0] data_out_7_lpi_3;
  reg [15:0] data_out_57_lpi_3;
  reg [15:0] data_out_5_lpi_3;
  reg [15:0] data_out_59_lpi_3;
  reg [15:0] data_out_3_lpi_3;
  reg [15:0] data_out_61_lpi_3;
  reg [15:0] data_out_1_lpi_3;
  reg [15:0] data_out_63_lpi_3;
  reg [5:0] LOOPJ1_j_sva;
  reg [1023:0] q_channel_data_sva;
  reg [37:0] maxn_sva;
  reg [37:0] sum_array_27_lpi_5;
  reg [37:0] sum_array_28_lpi_5;
  reg [37:0] sum_array_26_lpi_5;
  reg [37:0] sum_array_29_lpi_5;
  reg [37:0] sum_array_25_lpi_5;
  reg [37:0] sum_array_30_lpi_5;
  reg [37:0] sum_array_24_lpi_5;
  reg [37:0] sum_array_31_lpi_5;
  reg [37:0] sum_array_23_lpi_5;
  reg [37:0] sum_array_32_lpi_5;
  reg [37:0] sum_array_22_lpi_5;
  reg [37:0] sum_array_33_lpi_5;
  reg [37:0] sum_array_21_lpi_5;
  reg [37:0] sum_array_34_lpi_5;
  reg [37:0] sum_array_20_lpi_5;
  reg [37:0] sum_array_35_lpi_5;
  reg [37:0] sum_array_19_lpi_5;
  reg [37:0] sum_array_36_lpi_5;
  reg [37:0] sum_array_18_lpi_5;
  reg [37:0] sum_array_37_lpi_5;
  reg [37:0] sum_array_17_lpi_5;
  reg [37:0] sum_array_38_lpi_5;
  reg [37:0] sum_array_16_lpi_5;
  reg [37:0] sum_array_39_lpi_5;
  reg [37:0] sum_array_15_lpi_5;
  reg [37:0] sum_array_40_lpi_5;
  reg [37:0] sum_array_14_lpi_5;
  reg [37:0] sum_array_41_lpi_5;
  reg [37:0] sum_array_13_lpi_5;
  reg [37:0] sum_array_42_lpi_5;
  reg [37:0] sum_array_12_lpi_5;
  reg [37:0] sum_array_43_lpi_5;
  reg [37:0] sum_array_11_lpi_5;
  reg [37:0] sum_array_44_lpi_5;
  reg [37:0] sum_array_10_lpi_5;
  reg [37:0] sum_array_45_lpi_5;
  reg [37:0] sum_array_9_lpi_5;
  reg [37:0] sum_array_46_lpi_5;
  reg [37:0] sum_array_8_lpi_5;
  reg [37:0] sum_array_47_lpi_5;
  reg [37:0] sum_array_7_lpi_5;
  reg [37:0] sum_array_48_lpi_5;
  reg [37:0] sum_array_6_lpi_5;
  reg [37:0] sum_array_49_lpi_5;
  reg [37:0] sum_array_5_lpi_5;
  reg [37:0] sum_array_50_lpi_5;
  reg [37:0] sum_array_4_lpi_5;
  reg [37:0] sum_array_51_lpi_5;
  reg [37:0] sum_array_3_lpi_5;
  reg [37:0] sum_array_52_lpi_5;
  reg [37:0] sum_array_2_lpi_5;
  reg [37:0] sum_array_53_lpi_5;
  reg [37:0] sum_array_1_lpi_5;
  reg [37:0] sum_array_54_lpi_5;
  reg [37:0] sum_array_0_lpi_5;
  reg [37:0] sum_array_55_lpi_5;
  reg [1023:0] k_channel_data_sva;
  reg [37:0] LOOPL1_ac_int_cctor_sva;
  reg [15:0] LOOPJ1_sum2_1_sva;
  reg [15:0] data_out_0_lpi_6;
  wire [37:0] sum_array_55_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_0_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_54_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_1_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_53_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_2_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_52_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_3_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_51_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_4_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_50_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_5_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_49_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_6_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_48_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_7_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_47_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_8_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_46_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_9_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_45_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_10_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_44_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_11_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_43_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_12_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_42_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_13_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_41_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_14_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_40_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_15_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_39_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_16_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_38_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_17_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_37_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_18_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_36_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_19_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_35_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_20_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_34_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_21_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_33_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_22_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_32_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_23_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_31_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_24_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_30_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_25_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_29_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_26_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_28_lpi_5_dfm_1_mx0w1;
  wire [37:0] sum_array_27_lpi_5_dfm_1_mx0w1;
  wire LOOPK2_else_nor_tmp_1;
  wire LOOPK2_else_LOOPK2_else_and_cse_1;
  wire LOOPK2_else_LOOPK2_else_and_1_cse_1;
  wire LOOPK2_else_LOOPK2_else_and_2_cse_1;
  wire LOOPK2_else_LOOPK2_else_and_3_cse_1;
  wire LOOPK2_else_LOOPK2_else_and_4_cse_1;
  wire [37:0] LOOPK2_acc_ncse_sva_1;
  wire [38:0] nl_LOOPK2_acc_ncse_sva_1;
  wire [4:0] operator_4_false_acc_psp_sva_1;
  wire [5:0] nl_operator_4_false_acc_psp_sva_1;
  wire [37:0] LOOPK2_mux_169;
  wire LOOPK3_exs_66_0;
  wire LOOPK3_exs_68_0;
  wire LOOPK3_exs_70_0;
  wire LOOPK3_exs_72_0;
  wire LOOPK3_exs_74_0;
  wire LOOPK3_exs_76_0;
  wire LOOPK3_exs_78_0;
  wire LOOPK3_exs_80_0;
  wire LOOPK3_exs_82_0;
  wire LOOPK3_exs_84_0;
  wire LOOPK3_exs_86_0;
  wire LOOPK3_exs_88_0;
  wire LOOPK3_exs_90_0;
  wire LOOPK3_exs_92_0;
  wire LOOPK3_exs_94_0;
  wire LOOPK3_exs_96_0;
  wire LOOPK3_exs_98_0;
  wire LOOPK3_exs_100_0;
  wire LOOPK3_exs_102_0;
  wire LOOPK3_exs_104_0;
  wire LOOPK3_exs_106_0;
  wire LOOPK3_exs_108_0;
  wire LOOPK3_exs_110_0;
  wire LOOPK3_exs_112_0;
  wire LOOPK3_exs_114_0;
  wire LOOPK3_exs_116_0;
  wire LOOPK3_exs_118_0;
  wire LOOPK3_exs_120_0;
  wire LOOPK3_exs_122_0;
  wire LOOPK3_exs_124_0;
  wire LOOPK3_exs_126_0;
  wire and_1639_rgt;
  wire LOOPK1_and_61_cse;
  wire LOOPI1_i_or_cse;
  wire [5:0] LOOPK5_mux_cse;
  wire or_tmp_759;
  wire or_tmp_766;
  wire or_tmp_773;
  wire or_tmp_780;
  wire or_tmp_787;
  wire or_tmp_794;
  wire or_tmp_801;
  wire or_tmp_808;
  wire or_tmp_815;
  wire or_tmp_822;
  wire or_tmp_829;
  wire or_tmp_836;
  wire or_tmp_843;
  wire or_tmp_850;
  wire or_tmp_857;
  wire or_tmp_868;
  wire or_tmp_873;
  wire or_tmp_878;
  wire or_tmp_883;
  wire or_tmp_888;
  wire or_tmp_893;
  wire or_tmp_898;
  wire or_tmp_903;
  wire or_tmp_908;
  wire or_tmp_913;
  wire or_tmp_918;
  wire or_tmp_923;
  wire or_tmp_928;
  wire or_tmp_933;
  wire or_tmp_938;
  wire or_tmp_943;
  wire or_tmp_948;
  wire or_tmp_953;
  wire or_tmp_958;
  wire or_tmp_963;
  wire or_tmp_968;
  wire or_tmp_973;
  wire or_tmp_978;
  wire or_tmp_983;
  wire or_tmp_988;
  wire or_tmp_993;
  wire or_tmp_998;
  wire or_tmp_1003;
  wire or_tmp_1008;
  wire or_tmp_1012;
  wire LOOPK2_if_1_equal_1_tmp;
  wire not_tmp_714;
  wire mux_tmp_46;
  wire nand_34_cse;
  wire nand_47_cse;
  wire nand_58_cse;
  wire nand_75_cse;
  wire nand_84_cse;
  wire or_1735_cse;
  wire and_2169_cse;
  wire nor_178_cse;
  wire nor_177_cse;
  wire nor_240_cse;
  wire nor_169_cse;
  wire nand_55_cse;
  wire nand_22_cse;
  wire nor_14_cse;
  wire nand_31_cse;
  wire nand_44_cse;
  wire nor_174_cse;
  wire nand_108_cse;
  wire nand_117_cse;
  wire nand_122_cse;
  wire and_2155_cse;
  wire or_1253_itm;
  wire [15:0] LOOPL1_mux_1_itm;
  wire operator_38_true_acc_itm_36;

  wire[3:0] operator_4_false_acc_nl;
  wire[4:0] nl_operator_4_false_acc_nl;
  wire LOOPI1_i_not_1_nl;
  wire not_254_nl;
  wire and_675_nl;
  wire and_677_nl;
  wire and_679_nl;
  wire and_684_nl;
  wire and_686_nl;
  wire and_688_nl;
  wire and_693_nl;
  wire and_695_nl;
  wire and_697_nl;
  wire and_702_nl;
  wire and_704_nl;
  wire and_706_nl;
  wire and_711_nl;
  wire and_713_nl;
  wire and_715_nl;
  wire and_720_nl;
  wire and_722_nl;
  wire and_724_nl;
  wire and_729_nl;
  wire and_731_nl;
  wire and_733_nl;
  wire and_738_nl;
  wire and_740_nl;
  wire and_742_nl;
  wire and_747_nl;
  wire and_749_nl;
  wire and_751_nl;
  wire and_756_nl;
  wire and_758_nl;
  wire and_760_nl;
  wire and_765_nl;
  wire and_767_nl;
  wire and_769_nl;
  wire and_774_nl;
  wire and_776_nl;
  wire and_778_nl;
  wire and_783_nl;
  wire and_785_nl;
  wire and_787_nl;
  wire and_792_nl;
  wire and_794_nl;
  wire and_796_nl;
  wire and_801_nl;
  wire and_803_nl;
  wire and_805_nl;
  wire and_810_nl;
  wire and_812_nl;
  wire and_814_nl;
  wire and_819_nl;
  wire and_821_nl;
  wire and_823_nl;
  wire and_828_nl;
  wire and_830_nl;
  wire and_832_nl;
  wire and_837_nl;
  wire and_839_nl;
  wire and_841_nl;
  wire and_846_nl;
  wire and_848_nl;
  wire and_850_nl;
  wire and_855_nl;
  wire and_857_nl;
  wire and_859_nl;
  wire and_864_nl;
  wire and_866_nl;
  wire and_868_nl;
  wire and_873_nl;
  wire and_875_nl;
  wire and_877_nl;
  wire and_882_nl;
  wire and_884_nl;
  wire and_886_nl;
  wire and_891_nl;
  wire and_893_nl;
  wire and_895_nl;
  wire and_900_nl;
  wire and_902_nl;
  wire and_904_nl;
  wire and_909_nl;
  wire and_911_nl;
  wire and_913_nl;
  wire and_918_nl;
  wire and_920_nl;
  wire and_922_nl;
  wire and_927_nl;
  wire and_929_nl;
  wire and_931_nl;
  wire and_936_nl;
  wire and_938_nl;
  wire and_940_nl;
  wire and_945_nl;
  wire and_947_nl;
  wire and_949_nl;
  wire and_954_nl;
  wire and_956_nl;
  wire and_958_nl;
  wire and_963_nl;
  wire and_965_nl;
  wire and_967_nl;
  wire and_972_nl;
  wire and_974_nl;
  wire and_976_nl;
  wire and_981_nl;
  wire and_983_nl;
  wire and_985_nl;
  wire and_990_nl;
  wire and_992_nl;
  wire and_994_nl;
  wire and_999_nl;
  wire and_1001_nl;
  wire and_1003_nl;
  wire and_1008_nl;
  wire and_1010_nl;
  wire and_1012_nl;
  wire and_1017_nl;
  wire and_1019_nl;
  wire and_1021_nl;
  wire and_1026_nl;
  wire and_1028_nl;
  wire and_1030_nl;
  wire and_1035_nl;
  wire and_1037_nl;
  wire and_1039_nl;
  wire and_1044_nl;
  wire and_1046_nl;
  wire and_1048_nl;
  wire and_1053_nl;
  wire and_1055_nl;
  wire and_1057_nl;
  wire and_1062_nl;
  wire and_1064_nl;
  wire and_1066_nl;
  wire and_1071_nl;
  wire and_1073_nl;
  wire and_1075_nl;
  wire and_1080_nl;
  wire and_1082_nl;
  wire and_1084_nl;
  wire and_1089_nl;
  wire and_1091_nl;
  wire and_1093_nl;
  wire and_1098_nl;
  wire and_1100_nl;
  wire and_1102_nl;
  wire and_1107_nl;
  wire and_1109_nl;
  wire and_1111_nl;
  wire and_1116_nl;
  wire and_1118_nl;
  wire and_1120_nl;
  wire and_1125_nl;
  wire and_1127_nl;
  wire and_1129_nl;
  wire and_1134_nl;
  wire and_1136_nl;
  wire and_1138_nl;
  wire and_1143_nl;
  wire and_1145_nl;
  wire and_1147_nl;
  wire and_1152_nl;
  wire and_1154_nl;
  wire and_1156_nl;
  wire and_1161_nl;
  wire and_1163_nl;
  wire and_1165_nl;
  wire and_1170_nl;
  wire and_1172_nl;
  wire and_1174_nl;
  wire[15:0] LOOPK3_and_60_nl;
  wire and_1178_nl;
  wire mux_nl;
  wire nor_144_nl;
  wire or_nl;
  wire[15:0] LOOPK3_and_61_nl;
  wire and_1185_nl;
  wire[15:0] LOOPK3_and_62_nl;
  wire and_1192_nl;
  wire mux_6_nl;
  wire nor_145_nl;
  wire or_1275_nl;
  wire[15:0] LOOPK3_and_63_nl;
  wire and_1199_nl;
  wire[15:0] LOOPK3_and_64_nl;
  wire and_1206_nl;
  wire mux_7_nl;
  wire nor_146_nl;
  wire or_1282_nl;
  wire[15:0] LOOPK3_and_65_nl;
  wire and_1213_nl;
  wire[15:0] LOOPK3_and_66_nl;
  wire and_1220_nl;
  wire mux_8_nl;
  wire nor_147_nl;
  wire or_1289_nl;
  wire[15:0] LOOPK3_and_67_nl;
  wire and_1227_nl;
  wire[15:0] LOOPK3_and_68_nl;
  wire and_1234_nl;
  wire mux_9_nl;
  wire nor_148_nl;
  wire or_1296_nl;
  wire[15:0] LOOPK3_and_69_nl;
  wire and_1241_nl;
  wire[15:0] LOOPK3_and_70_nl;
  wire and_1248_nl;
  wire mux_10_nl;
  wire nor_149_nl;
  wire or_1303_nl;
  wire[15:0] LOOPK3_and_71_nl;
  wire and_1255_nl;
  wire[15:0] LOOPK3_and_72_nl;
  wire and_1262_nl;
  wire mux_11_nl;
  wire nor_150_nl;
  wire or_1310_nl;
  wire[15:0] LOOPK3_and_73_nl;
  wire and_1269_nl;
  wire[15:0] LOOPK3_and_74_nl;
  wire and_1276_nl;
  wire mux_12_nl;
  wire nor_151_nl;
  wire[15:0] LOOPK3_and_75_nl;
  wire and_1283_nl;
  wire[15:0] LOOPK3_and_76_nl;
  wire and_1290_nl;
  wire mux_13_nl;
  wire and_2736_nl;
  wire or_1324_nl;
  wire[15:0] LOOPK3_and_77_nl;
  wire and_1297_nl;
  wire[15:0] LOOPK3_and_78_nl;
  wire and_1304_nl;
  wire mux_14_nl;
  wire and_2738_nl;
  wire or_1331_nl;
  wire[15:0] LOOPK3_and_79_nl;
  wire and_1311_nl;
  wire[15:0] LOOPK3_and_80_nl;
  wire and_1318_nl;
  wire mux_15_nl;
  wire and_2740_nl;
  wire or_1338_nl;
  wire[15:0] LOOPK3_and_81_nl;
  wire and_1325_nl;
  wire[15:0] LOOPK3_and_82_nl;
  wire and_1332_nl;
  wire mux_16_nl;
  wire and_2742_nl;
  wire[15:0] LOOPK3_and_83_nl;
  wire and_1339_nl;
  wire[15:0] LOOPK3_and_84_nl;
  wire and_1346_nl;
  wire mux_17_nl;
  wire and_2744_nl;
  wire or_1352_nl;
  wire[15:0] LOOPK3_and_85_nl;
  wire and_1353_nl;
  wire[15:0] LOOPK3_and_86_nl;
  wire and_1360_nl;
  wire mux_18_nl;
  wire and_2746_nl;
  wire or_1359_nl;
  wire[15:0] LOOPK3_and_87_nl;
  wire and_1367_nl;
  wire[15:0] LOOPK3_and_88_nl;
  wire and_1374_nl;
  wire mux_19_nl;
  wire and_2748_nl;
  wire or_1366_nl;
  wire[15:0] LOOPK3_and_89_nl;
  wire and_1381_nl;
  wire[15:0] LOOPK3_and_90_nl;
  wire and_1388_nl;
  wire[15:0] LOOPK3_and_152_nl;
  wire and_1395_nl;
  wire mux_20_nl;
  wire nor_153_nl;
  wire nand_56_nl;
  wire[15:0] LOOPK3_and_153_nl;
  wire and_1402_nl;
  wire mux_21_nl;
  wire and_2752_nl;
  wire or_1381_nl;
  wire[15:0] LOOPK3_and_154_nl;
  wire and_1409_nl;
  wire mux_22_nl;
  wire nor_154_nl;
  wire or_1386_nl;
  wire[15:0] LOOPK3_and_155_nl;
  wire and_1416_nl;
  wire mux_23_nl;
  wire and_2754_nl;
  wire or_1391_nl;
  wire[15:0] LOOPK3_and_156_nl;
  wire and_1423_nl;
  wire mux_24_nl;
  wire nor_155_nl;
  wire or_1396_nl;
  wire[15:0] LOOPK3_and_157_nl;
  wire and_1430_nl;
  wire mux_25_nl;
  wire and_2756_nl;
  wire or_1401_nl;
  wire[15:0] LOOPK3_and_158_nl;
  wire and_1437_nl;
  wire mux_26_nl;
  wire nor_156_nl;
  wire or_1406_nl;
  wire[15:0] LOOPK3_and_159_nl;
  wire and_1444_nl;
  wire mux_27_nl;
  wire and_2758_nl;
  wire or_1411_nl;
  wire[15:0] LOOPK3_and_160_nl;
  wire and_1451_nl;
  wire mux_28_nl;
  wire nor_157_nl;
  wire or_1416_nl;
  wire[15:0] LOOPK3_and_161_nl;
  wire and_1458_nl;
  wire mux_29_nl;
  wire and_2760_nl;
  wire or_1421_nl;
  wire[15:0] LOOPK3_and_162_nl;
  wire and_1465_nl;
  wire mux_30_nl;
  wire nor_158_nl;
  wire or_1426_nl;
  wire[15:0] LOOPK3_and_163_nl;
  wire and_1472_nl;
  wire mux_31_nl;
  wire and_2762_nl;
  wire or_1431_nl;
  wire[15:0] LOOPK3_and_164_nl;
  wire and_1479_nl;
  wire mux_32_nl;
  wire nor_159_nl;
  wire or_1436_nl;
  wire[15:0] LOOPK3_and_165_nl;
  wire and_1486_nl;
  wire mux_33_nl;
  wire and_2764_nl;
  wire or_1441_nl;
  wire[15:0] LOOPK3_and_166_nl;
  wire and_1493_nl;
  wire mux_34_nl;
  wire nor_160_nl;
  wire or_1446_nl;
  wire[15:0] LOOPK3_and_167_nl;
  wire and_1500_nl;
  wire mux_35_nl;
  wire and_2766_nl;
  wire nand_73_nl;
  wire[15:0] LOOPK3_and_168_nl;
  wire and_1507_nl;
  wire mux_36_nl;
  wire nor_161_nl;
  wire or_1456_nl;
  wire[15:0] LOOPK3_and_169_nl;
  wire and_1514_nl;
  wire mux_37_nl;
  wire and_2768_nl;
  wire or_1461_nl;
  wire[15:0] LOOPK3_and_170_nl;
  wire and_1521_nl;
  wire mux_38_nl;
  wire nor_162_nl;
  wire or_1466_nl;
  wire[15:0] LOOPK3_and_171_nl;
  wire and_1528_nl;
  wire mux_39_nl;
  wire and_2770_nl;
  wire or_1471_nl;
  wire[15:0] LOOPK3_and_172_nl;
  wire and_1535_nl;
  wire mux_40_nl;
  wire nor_163_nl;
  wire or_1476_nl;
  wire[15:0] LOOPK3_and_173_nl;
  wire and_1542_nl;
  wire mux_41_nl;
  wire and_2772_nl;
  wire or_1481_nl;
  wire[15:0] LOOPK3_and_174_nl;
  wire and_1549_nl;
  wire mux_42_nl;
  wire nor_164_nl;
  wire or_1486_nl;
  wire[15:0] LOOPK3_and_175_nl;
  wire and_1556_nl;
  wire mux_43_nl;
  wire and_2774_nl;
  wire nand_82_nl;
  wire[15:0] LOOPK3_and_176_nl;
  wire and_1563_nl;
  wire mux_44_nl;
  wire nor_165_nl;
  wire or_1496_nl;
  wire[15:0] LOOPK3_and_177_nl;
  wire and_1570_nl;
  wire mux_45_nl;
  wire and_2776_nl;
  wire or_1501_nl;
  wire[15:0] LOOPK3_and_178_nl;
  wire and_1577_nl;
  wire mux_46_nl;
  wire nor_166_nl;
  wire or_1506_nl;
  wire[15:0] LOOPK3_and_179_nl;
  wire and_1584_nl;
  wire mux_47_nl;
  wire and_2778_nl;
  wire or_1511_nl;
  wire[15:0] LOOPK3_and_180_nl;
  wire and_1591_nl;
  wire mux_48_nl;
  wire nor_167_nl;
  wire or_1516_nl;
  wire[15:0] LOOPK3_and_181_nl;
  wire and_1598_nl;
  wire mux_49_nl;
  wire and_2780_nl;
  wire[15:0] nor_402_nl;
  wire data_out_or_63_nl;
  wire or_1744_nl;
  wire[15:0] LOOPK3_and_183_nl;
  wire and_1614_nl;
  wire cnt_nor_nl;
  wire[38:0] LOOPK1_acc_1_nl;
  wire[39:0] nl_LOOPK1_acc_1_nl;
  wire LOOPK1_endflag_mux1h_2_nl;
  wire LOOPK3_if_LOOPK3_if_and_nl;
  wire LOOPL1_l_LOOPL1_l_mux_nl;
  wire[5:0] LOOPL1_l_LOOPL1_l_mux_1_nl;
  wire or_1232_nl;
  wire and_2822_nl;
  wire mux_52_nl;
  wire mux_51_nl;
  wire or_1732_nl;
  wire or_1736_nl;
  wire[37:0] LOOPL1_acc_nl;
  wire[38:0] nl_LOOPL1_acc_nl;
  wire[15:0] LOOPJ1_sum2_mux_nl;
  wire[15:0] operator_16_false_div_nl;
  wire not_370_nl;
  wire data_out_nand_nl;
  wire[31:0] LOOPL2_acc_1_nl;
  wire[32:0] nl_LOOPL2_acc_1_nl;
  wire[37:0] LOOPK2_if_and_171_nl;
  wire LOOPK2_if_not_232_nl;
  wire LOOPK2_LOOPK2_nor_56_nl;
  wire LOOPK2_else_and_1981_nl;
  wire LOOPK2_else_and_1983_nl;
  wire LOOPK2_else_and_1985_nl;
  wire LOOPK2_else_and_1987_nl;
  wire LOOPK2_else_and_1989_nl;
  wire LOOPK2_else_and_1991_nl;
  wire LOOPK2_else_and_1993_nl;
  wire LOOPK2_else_and_1995_nl;
  wire LOOPK2_else_and_1997_nl;
  wire LOOPK2_else_and_1999_nl;
  wire LOOPK2_else_and_2001_nl;
  wire LOOPK2_else_and_2003_nl;
  wire LOOPK2_else_and_2005_nl;
  wire LOOPK2_else_and_2007_nl;
  wire LOOPK2_else_and_2009_nl;
  wire LOOPK2_else_and_2011_nl;
  wire LOOPK2_else_and_2013_nl;
  wire LOOPK2_else_and_2015_nl;
  wire[37:0] LOOPK2_if_and_170_nl;
  wire LOOPK2_if_not_250_nl;
  wire LOOPK2_LOOPK2_nor_1_nl;
  wire LOOPK2_else_and_1_nl;
  wire LOOPK2_else_and_3_nl;
  wire LOOPK2_else_and_5_nl;
  wire LOOPK2_else_and_7_nl;
  wire LOOPK2_else_and_9_nl;
  wire LOOPK2_else_and_11_nl;
  wire LOOPK2_else_and_13_nl;
  wire LOOPK2_else_and_15_nl;
  wire LOOPK2_else_and_17_nl;
  wire LOOPK2_else_and_19_nl;
  wire LOOPK2_else_and_21_nl;
  wire LOOPK2_else_and_23_nl;
  wire LOOPK2_else_and_25_nl;
  wire LOOPK2_else_and_27_nl;
  wire LOOPK2_else_and_29_nl;
  wire LOOPK2_else_and_31_nl;
  wire LOOPK2_else_and_33_nl;
  wire LOOPK2_else_and_35_nl;
  wire[37:0] LOOPK2_if_and_169_nl;
  wire LOOPK2_if_not_268_nl;
  wire LOOPK2_LOOPK2_nor_55_nl;
  wire LOOPK2_else_and_1945_nl;
  wire LOOPK2_else_and_1947_nl;
  wire LOOPK2_else_and_1949_nl;
  wire LOOPK2_else_and_1951_nl;
  wire LOOPK2_else_and_1953_nl;
  wire LOOPK2_else_and_1955_nl;
  wire LOOPK2_else_and_1957_nl;
  wire LOOPK2_else_and_1959_nl;
  wire LOOPK2_else_and_1961_nl;
  wire LOOPK2_else_and_1963_nl;
  wire LOOPK2_else_and_1965_nl;
  wire LOOPK2_else_and_1967_nl;
  wire LOOPK2_else_and_1969_nl;
  wire LOOPK2_else_and_1971_nl;
  wire LOOPK2_else_and_1973_nl;
  wire LOOPK2_else_and_1975_nl;
  wire LOOPK2_else_and_1977_nl;
  wire LOOPK2_else_and_1979_nl;
  wire[37:0] LOOPK2_if_and_168_nl;
  wire LOOPK2_if_not_286_nl;
  wire LOOPK2_LOOPK2_nor_2_nl;
  wire LOOPK2_else_and_37_nl;
  wire LOOPK2_else_and_39_nl;
  wire LOOPK2_else_and_41_nl;
  wire LOOPK2_else_and_43_nl;
  wire LOOPK2_else_and_45_nl;
  wire LOOPK2_else_and_47_nl;
  wire LOOPK2_else_and_49_nl;
  wire LOOPK2_else_and_51_nl;
  wire LOOPK2_else_and_53_nl;
  wire LOOPK2_else_and_55_nl;
  wire LOOPK2_else_and_57_nl;
  wire LOOPK2_else_and_59_nl;
  wire LOOPK2_else_and_61_nl;
  wire LOOPK2_else_and_63_nl;
  wire LOOPK2_else_and_65_nl;
  wire LOOPK2_else_and_67_nl;
  wire LOOPK2_else_and_69_nl;
  wire LOOPK2_else_and_71_nl;
  wire[37:0] LOOPK2_if_and_167_nl;
  wire LOOPK2_if_not_304_nl;
  wire LOOPK2_LOOPK2_nor_54_nl;
  wire LOOPK2_else_and_1909_nl;
  wire LOOPK2_else_and_1911_nl;
  wire LOOPK2_else_and_1913_nl;
  wire LOOPK2_else_and_1915_nl;
  wire LOOPK2_else_and_1917_nl;
  wire LOOPK2_else_and_1919_nl;
  wire LOOPK2_else_and_1921_nl;
  wire LOOPK2_else_and_1923_nl;
  wire LOOPK2_else_and_1925_nl;
  wire LOOPK2_else_and_1927_nl;
  wire LOOPK2_else_and_1929_nl;
  wire LOOPK2_else_and_1931_nl;
  wire LOOPK2_else_and_1933_nl;
  wire LOOPK2_else_and_1935_nl;
  wire LOOPK2_else_and_1937_nl;
  wire LOOPK2_else_and_1939_nl;
  wire LOOPK2_else_and_1941_nl;
  wire LOOPK2_else_and_1943_nl;
  wire[37:0] LOOPK2_if_and_166_nl;
  wire LOOPK2_if_not_322_nl;
  wire LOOPK2_LOOPK2_nor_3_nl;
  wire LOOPK2_else_and_73_nl;
  wire LOOPK2_else_and_75_nl;
  wire LOOPK2_else_and_77_nl;
  wire LOOPK2_else_and_79_nl;
  wire LOOPK2_else_and_81_nl;
  wire LOOPK2_else_and_83_nl;
  wire LOOPK2_else_and_85_nl;
  wire LOOPK2_else_and_87_nl;
  wire LOOPK2_else_and_89_nl;
  wire LOOPK2_else_and_91_nl;
  wire LOOPK2_else_and_93_nl;
  wire LOOPK2_else_and_95_nl;
  wire LOOPK2_else_and_97_nl;
  wire LOOPK2_else_and_99_nl;
  wire LOOPK2_else_and_101_nl;
  wire LOOPK2_else_and_103_nl;
  wire LOOPK2_else_and_105_nl;
  wire LOOPK2_else_and_107_nl;
  wire[37:0] LOOPK2_if_and_165_nl;
  wire LOOPK2_if_not_340_nl;
  wire LOOPK2_LOOPK2_nor_53_nl;
  wire LOOPK2_else_and_1873_nl;
  wire LOOPK2_else_and_1875_nl;
  wire LOOPK2_else_and_1877_nl;
  wire LOOPK2_else_and_1879_nl;
  wire LOOPK2_else_and_1881_nl;
  wire LOOPK2_else_and_1883_nl;
  wire LOOPK2_else_and_1885_nl;
  wire LOOPK2_else_and_1887_nl;
  wire LOOPK2_else_and_1889_nl;
  wire LOOPK2_else_and_1891_nl;
  wire LOOPK2_else_and_1893_nl;
  wire LOOPK2_else_and_1895_nl;
  wire LOOPK2_else_and_1897_nl;
  wire LOOPK2_else_and_1899_nl;
  wire LOOPK2_else_and_1901_nl;
  wire LOOPK2_else_and_1903_nl;
  wire LOOPK2_else_and_1905_nl;
  wire LOOPK2_else_and_1907_nl;
  wire[37:0] LOOPK2_if_and_164_nl;
  wire LOOPK2_if_not_358_nl;
  wire LOOPK2_LOOPK2_nor_4_nl;
  wire LOOPK2_else_and_109_nl;
  wire LOOPK2_else_and_111_nl;
  wire LOOPK2_else_and_113_nl;
  wire LOOPK2_else_and_115_nl;
  wire LOOPK2_else_and_117_nl;
  wire LOOPK2_else_and_119_nl;
  wire LOOPK2_else_and_121_nl;
  wire LOOPK2_else_and_123_nl;
  wire LOOPK2_else_and_125_nl;
  wire LOOPK2_else_and_127_nl;
  wire LOOPK2_else_and_129_nl;
  wire LOOPK2_else_and_131_nl;
  wire LOOPK2_else_and_133_nl;
  wire LOOPK2_else_and_135_nl;
  wire LOOPK2_else_and_137_nl;
  wire LOOPK2_else_and_139_nl;
  wire LOOPK2_else_and_141_nl;
  wire LOOPK2_else_and_143_nl;
  wire[37:0] LOOPK2_if_and_163_nl;
  wire LOOPK2_if_not_376_nl;
  wire LOOPK2_LOOPK2_nor_52_nl;
  wire LOOPK2_else_and_1837_nl;
  wire LOOPK2_else_and_1839_nl;
  wire LOOPK2_else_and_1841_nl;
  wire LOOPK2_else_and_1843_nl;
  wire LOOPK2_else_and_1845_nl;
  wire LOOPK2_else_and_1847_nl;
  wire LOOPK2_else_and_1849_nl;
  wire LOOPK2_else_and_1851_nl;
  wire LOOPK2_else_and_1853_nl;
  wire LOOPK2_else_and_1855_nl;
  wire LOOPK2_else_and_1857_nl;
  wire LOOPK2_else_and_1859_nl;
  wire LOOPK2_else_and_1861_nl;
  wire LOOPK2_else_and_1863_nl;
  wire LOOPK2_else_and_1865_nl;
  wire LOOPK2_else_and_1867_nl;
  wire LOOPK2_else_and_1869_nl;
  wire LOOPK2_else_and_1871_nl;
  wire[37:0] LOOPK2_if_and_162_nl;
  wire LOOPK2_if_not_394_nl;
  wire LOOPK2_LOOPK2_nor_5_nl;
  wire LOOPK2_else_and_145_nl;
  wire LOOPK2_else_and_147_nl;
  wire LOOPK2_else_and_149_nl;
  wire LOOPK2_else_and_151_nl;
  wire LOOPK2_else_and_153_nl;
  wire LOOPK2_else_and_155_nl;
  wire LOOPK2_else_and_157_nl;
  wire LOOPK2_else_and_159_nl;
  wire LOOPK2_else_and_161_nl;
  wire LOOPK2_else_and_163_nl;
  wire LOOPK2_else_and_165_nl;
  wire LOOPK2_else_and_167_nl;
  wire LOOPK2_else_and_169_nl;
  wire LOOPK2_else_and_171_nl;
  wire LOOPK2_else_and_173_nl;
  wire LOOPK2_else_and_175_nl;
  wire LOOPK2_else_and_177_nl;
  wire LOOPK2_else_and_179_nl;
  wire[37:0] LOOPK2_if_and_161_nl;
  wire LOOPK2_if_not_412_nl;
  wire LOOPK2_LOOPK2_nor_51_nl;
  wire LOOPK2_else_and_1801_nl;
  wire LOOPK2_else_and_1803_nl;
  wire LOOPK2_else_and_1805_nl;
  wire LOOPK2_else_and_1807_nl;
  wire LOOPK2_else_and_1809_nl;
  wire LOOPK2_else_and_1811_nl;
  wire LOOPK2_else_and_1813_nl;
  wire LOOPK2_else_and_1815_nl;
  wire LOOPK2_else_and_1817_nl;
  wire LOOPK2_else_and_1819_nl;
  wire LOOPK2_else_and_1821_nl;
  wire LOOPK2_else_and_1823_nl;
  wire LOOPK2_else_and_1825_nl;
  wire LOOPK2_else_and_1827_nl;
  wire LOOPK2_else_and_1829_nl;
  wire LOOPK2_else_and_1831_nl;
  wire LOOPK2_else_and_1833_nl;
  wire LOOPK2_else_and_1835_nl;
  wire[37:0] LOOPK2_if_and_160_nl;
  wire LOOPK2_if_not_430_nl;
  wire LOOPK2_LOOPK2_nor_6_nl;
  wire LOOPK2_else_and_181_nl;
  wire LOOPK2_else_and_183_nl;
  wire LOOPK2_else_and_185_nl;
  wire LOOPK2_else_and_187_nl;
  wire LOOPK2_else_and_189_nl;
  wire LOOPK2_else_and_191_nl;
  wire LOOPK2_else_and_193_nl;
  wire LOOPK2_else_and_195_nl;
  wire LOOPK2_else_and_197_nl;
  wire LOOPK2_else_and_199_nl;
  wire LOOPK2_else_and_201_nl;
  wire LOOPK2_else_and_203_nl;
  wire LOOPK2_else_and_205_nl;
  wire LOOPK2_else_and_207_nl;
  wire LOOPK2_else_and_209_nl;
  wire LOOPK2_else_and_211_nl;
  wire LOOPK2_else_and_213_nl;
  wire LOOPK2_else_and_215_nl;
  wire[37:0] LOOPK2_if_and_159_nl;
  wire LOOPK2_if_not_448_nl;
  wire LOOPK2_LOOPK2_nor_50_nl;
  wire LOOPK2_else_and_1765_nl;
  wire LOOPK2_else_and_1767_nl;
  wire LOOPK2_else_and_1769_nl;
  wire LOOPK2_else_and_1771_nl;
  wire LOOPK2_else_and_1773_nl;
  wire LOOPK2_else_and_1775_nl;
  wire LOOPK2_else_and_1777_nl;
  wire LOOPK2_else_and_1779_nl;
  wire LOOPK2_else_and_1781_nl;
  wire LOOPK2_else_and_1783_nl;
  wire LOOPK2_else_and_1785_nl;
  wire LOOPK2_else_and_1787_nl;
  wire LOOPK2_else_and_1789_nl;
  wire LOOPK2_else_and_1791_nl;
  wire LOOPK2_else_and_1793_nl;
  wire LOOPK2_else_and_1795_nl;
  wire LOOPK2_else_and_1797_nl;
  wire LOOPK2_else_and_1799_nl;
  wire[37:0] LOOPK2_if_and_158_nl;
  wire LOOPK2_if_not_466_nl;
  wire LOOPK2_LOOPK2_nor_7_nl;
  wire LOOPK2_else_and_217_nl;
  wire LOOPK2_else_and_219_nl;
  wire LOOPK2_else_and_221_nl;
  wire LOOPK2_else_and_223_nl;
  wire LOOPK2_else_and_225_nl;
  wire LOOPK2_else_and_227_nl;
  wire LOOPK2_else_and_229_nl;
  wire LOOPK2_else_and_231_nl;
  wire LOOPK2_else_and_233_nl;
  wire LOOPK2_else_and_235_nl;
  wire LOOPK2_else_and_237_nl;
  wire LOOPK2_else_and_239_nl;
  wire LOOPK2_else_and_241_nl;
  wire LOOPK2_else_and_243_nl;
  wire LOOPK2_else_and_245_nl;
  wire LOOPK2_else_and_247_nl;
  wire LOOPK2_else_and_249_nl;
  wire LOOPK2_else_and_251_nl;
  wire[37:0] LOOPK2_if_and_157_nl;
  wire LOOPK2_if_not_484_nl;
  wire LOOPK2_LOOPK2_nor_49_nl;
  wire LOOPK2_else_and_1729_nl;
  wire LOOPK2_else_and_1731_nl;
  wire LOOPK2_else_and_1733_nl;
  wire LOOPK2_else_and_1735_nl;
  wire LOOPK2_else_and_1737_nl;
  wire LOOPK2_else_and_1739_nl;
  wire LOOPK2_else_and_1741_nl;
  wire LOOPK2_else_and_1743_nl;
  wire LOOPK2_else_and_1745_nl;
  wire LOOPK2_else_and_1747_nl;
  wire LOOPK2_else_and_1749_nl;
  wire LOOPK2_else_and_1751_nl;
  wire LOOPK2_else_and_1753_nl;
  wire LOOPK2_else_and_1755_nl;
  wire LOOPK2_else_and_1757_nl;
  wire LOOPK2_else_and_1759_nl;
  wire LOOPK2_else_and_1761_nl;
  wire LOOPK2_else_and_1763_nl;
  wire[37:0] LOOPK2_if_and_156_nl;
  wire LOOPK2_if_not_502_nl;
  wire LOOPK2_LOOPK2_nor_8_nl;
  wire LOOPK2_else_and_253_nl;
  wire LOOPK2_else_and_255_nl;
  wire LOOPK2_else_and_257_nl;
  wire LOOPK2_else_and_259_nl;
  wire LOOPK2_else_and_261_nl;
  wire LOOPK2_else_and_263_nl;
  wire LOOPK2_else_and_265_nl;
  wire LOOPK2_else_and_267_nl;
  wire LOOPK2_else_and_269_nl;
  wire LOOPK2_else_and_271_nl;
  wire LOOPK2_else_and_273_nl;
  wire LOOPK2_else_and_275_nl;
  wire LOOPK2_else_and_277_nl;
  wire LOOPK2_else_and_279_nl;
  wire LOOPK2_else_and_281_nl;
  wire LOOPK2_else_and_283_nl;
  wire LOOPK2_else_and_285_nl;
  wire LOOPK2_else_and_287_nl;
  wire[37:0] LOOPK2_if_and_155_nl;
  wire LOOPK2_if_not_520_nl;
  wire LOOPK2_LOOPK2_nor_48_nl;
  wire LOOPK2_else_and_1693_nl;
  wire LOOPK2_else_and_1695_nl;
  wire LOOPK2_else_and_1697_nl;
  wire LOOPK2_else_and_1699_nl;
  wire LOOPK2_else_and_1701_nl;
  wire LOOPK2_else_and_1703_nl;
  wire LOOPK2_else_and_1705_nl;
  wire LOOPK2_else_and_1707_nl;
  wire LOOPK2_else_and_1709_nl;
  wire LOOPK2_else_and_1711_nl;
  wire LOOPK2_else_and_1713_nl;
  wire LOOPK2_else_and_1715_nl;
  wire LOOPK2_else_and_1717_nl;
  wire LOOPK2_else_and_1719_nl;
  wire LOOPK2_else_and_1721_nl;
  wire LOOPK2_else_and_1723_nl;
  wire LOOPK2_else_and_1725_nl;
  wire LOOPK2_else_and_1727_nl;
  wire[37:0] LOOPK2_if_and_154_nl;
  wire LOOPK2_if_not_538_nl;
  wire LOOPK2_LOOPK2_nor_9_nl;
  wire LOOPK2_else_and_289_nl;
  wire LOOPK2_else_and_291_nl;
  wire LOOPK2_else_and_293_nl;
  wire LOOPK2_else_and_295_nl;
  wire LOOPK2_else_and_297_nl;
  wire LOOPK2_else_and_299_nl;
  wire LOOPK2_else_and_301_nl;
  wire LOOPK2_else_and_303_nl;
  wire LOOPK2_else_and_305_nl;
  wire LOOPK2_else_and_307_nl;
  wire LOOPK2_else_and_309_nl;
  wire LOOPK2_else_and_311_nl;
  wire LOOPK2_else_and_313_nl;
  wire LOOPK2_else_and_315_nl;
  wire LOOPK2_else_and_317_nl;
  wire LOOPK2_else_and_319_nl;
  wire LOOPK2_else_and_321_nl;
  wire LOOPK2_else_and_323_nl;
  wire[37:0] LOOPK2_if_and_153_nl;
  wire LOOPK2_if_not_556_nl;
  wire LOOPK2_LOOPK2_nor_47_nl;
  wire LOOPK2_else_and_1657_nl;
  wire LOOPK2_else_and_1659_nl;
  wire LOOPK2_else_and_1661_nl;
  wire LOOPK2_else_and_1663_nl;
  wire LOOPK2_else_and_1665_nl;
  wire LOOPK2_else_and_1667_nl;
  wire LOOPK2_else_and_1669_nl;
  wire LOOPK2_else_and_1671_nl;
  wire LOOPK2_else_and_1673_nl;
  wire LOOPK2_else_and_1675_nl;
  wire LOOPK2_else_and_1677_nl;
  wire LOOPK2_else_and_1679_nl;
  wire LOOPK2_else_and_1681_nl;
  wire LOOPK2_else_and_1683_nl;
  wire LOOPK2_else_and_1685_nl;
  wire LOOPK2_else_and_1687_nl;
  wire LOOPK2_else_and_1689_nl;
  wire LOOPK2_else_and_1691_nl;
  wire[37:0] LOOPK2_if_and_152_nl;
  wire LOOPK2_if_not_574_nl;
  wire LOOPK2_LOOPK2_nor_10_nl;
  wire LOOPK2_else_and_325_nl;
  wire LOOPK2_else_and_327_nl;
  wire LOOPK2_else_and_329_nl;
  wire LOOPK2_else_and_331_nl;
  wire LOOPK2_else_and_333_nl;
  wire LOOPK2_else_and_335_nl;
  wire LOOPK2_else_and_337_nl;
  wire LOOPK2_else_and_339_nl;
  wire LOOPK2_else_and_341_nl;
  wire LOOPK2_else_and_343_nl;
  wire LOOPK2_else_and_345_nl;
  wire LOOPK2_else_and_347_nl;
  wire LOOPK2_else_and_349_nl;
  wire LOOPK2_else_and_351_nl;
  wire LOOPK2_else_and_353_nl;
  wire LOOPK2_else_and_355_nl;
  wire LOOPK2_else_and_357_nl;
  wire LOOPK2_else_and_359_nl;
  wire[37:0] LOOPK2_if_and_151_nl;
  wire LOOPK2_if_not_592_nl;
  wire LOOPK2_LOOPK2_nor_46_nl;
  wire LOOPK2_else_and_1621_nl;
  wire LOOPK2_else_and_1623_nl;
  wire LOOPK2_else_and_1625_nl;
  wire LOOPK2_else_and_1627_nl;
  wire LOOPK2_else_and_1629_nl;
  wire LOOPK2_else_and_1631_nl;
  wire LOOPK2_else_and_1633_nl;
  wire LOOPK2_else_and_1635_nl;
  wire LOOPK2_else_and_1637_nl;
  wire LOOPK2_else_and_1639_nl;
  wire LOOPK2_else_and_1641_nl;
  wire LOOPK2_else_and_1643_nl;
  wire LOOPK2_else_and_1645_nl;
  wire LOOPK2_else_and_1647_nl;
  wire LOOPK2_else_and_1649_nl;
  wire LOOPK2_else_and_1651_nl;
  wire LOOPK2_else_and_1653_nl;
  wire LOOPK2_else_and_1655_nl;
  wire[37:0] LOOPK2_if_and_150_nl;
  wire LOOPK2_if_not_610_nl;
  wire LOOPK2_LOOPK2_nor_11_nl;
  wire LOOPK2_else_and_361_nl;
  wire LOOPK2_else_and_363_nl;
  wire LOOPK2_else_and_365_nl;
  wire LOOPK2_else_and_367_nl;
  wire LOOPK2_else_and_369_nl;
  wire LOOPK2_else_and_371_nl;
  wire LOOPK2_else_and_373_nl;
  wire LOOPK2_else_and_375_nl;
  wire LOOPK2_else_and_377_nl;
  wire LOOPK2_else_and_379_nl;
  wire LOOPK2_else_and_381_nl;
  wire LOOPK2_else_and_383_nl;
  wire LOOPK2_else_and_385_nl;
  wire LOOPK2_else_and_387_nl;
  wire LOOPK2_else_and_389_nl;
  wire LOOPK2_else_and_391_nl;
  wire LOOPK2_else_and_393_nl;
  wire LOOPK2_else_and_395_nl;
  wire[37:0] LOOPK2_if_and_149_nl;
  wire LOOPK2_if_not_628_nl;
  wire LOOPK2_LOOPK2_nor_45_nl;
  wire LOOPK2_else_and_1585_nl;
  wire LOOPK2_else_and_1587_nl;
  wire LOOPK2_else_and_1589_nl;
  wire LOOPK2_else_and_1591_nl;
  wire LOOPK2_else_and_1593_nl;
  wire LOOPK2_else_and_1595_nl;
  wire LOOPK2_else_and_1597_nl;
  wire LOOPK2_else_and_1599_nl;
  wire LOOPK2_else_and_1601_nl;
  wire LOOPK2_else_and_1603_nl;
  wire LOOPK2_else_and_1605_nl;
  wire LOOPK2_else_and_1607_nl;
  wire LOOPK2_else_and_1609_nl;
  wire LOOPK2_else_and_1611_nl;
  wire LOOPK2_else_and_1613_nl;
  wire LOOPK2_else_and_1615_nl;
  wire LOOPK2_else_and_1617_nl;
  wire LOOPK2_else_and_1619_nl;
  wire[37:0] LOOPK2_if_and_148_nl;
  wire LOOPK2_if_not_646_nl;
  wire LOOPK2_LOOPK2_nor_12_nl;
  wire LOOPK2_else_and_397_nl;
  wire LOOPK2_else_and_399_nl;
  wire LOOPK2_else_and_401_nl;
  wire LOOPK2_else_and_403_nl;
  wire LOOPK2_else_and_405_nl;
  wire LOOPK2_else_and_407_nl;
  wire LOOPK2_else_and_409_nl;
  wire LOOPK2_else_and_411_nl;
  wire LOOPK2_else_and_413_nl;
  wire LOOPK2_else_and_415_nl;
  wire LOOPK2_else_and_417_nl;
  wire LOOPK2_else_and_419_nl;
  wire LOOPK2_else_and_421_nl;
  wire LOOPK2_else_and_423_nl;
  wire LOOPK2_else_and_425_nl;
  wire LOOPK2_else_and_427_nl;
  wire LOOPK2_else_and_429_nl;
  wire LOOPK2_else_and_431_nl;
  wire[37:0] LOOPK2_if_and_147_nl;
  wire LOOPK2_if_not_664_nl;
  wire LOOPK2_LOOPK2_nor_44_nl;
  wire LOOPK2_else_and_1549_nl;
  wire LOOPK2_else_and_1551_nl;
  wire LOOPK2_else_and_1553_nl;
  wire LOOPK2_else_and_1555_nl;
  wire LOOPK2_else_and_1557_nl;
  wire LOOPK2_else_and_1559_nl;
  wire LOOPK2_else_and_1561_nl;
  wire LOOPK2_else_and_1563_nl;
  wire LOOPK2_else_and_1565_nl;
  wire LOOPK2_else_and_1567_nl;
  wire LOOPK2_else_and_1569_nl;
  wire LOOPK2_else_and_1571_nl;
  wire LOOPK2_else_and_1573_nl;
  wire LOOPK2_else_and_1575_nl;
  wire LOOPK2_else_and_1577_nl;
  wire LOOPK2_else_and_1579_nl;
  wire LOOPK2_else_and_1581_nl;
  wire LOOPK2_else_and_1583_nl;
  wire[37:0] LOOPK2_if_and_146_nl;
  wire LOOPK2_if_not_682_nl;
  wire LOOPK2_LOOPK2_nor_13_nl;
  wire LOOPK2_else_and_433_nl;
  wire LOOPK2_else_and_435_nl;
  wire LOOPK2_else_and_437_nl;
  wire LOOPK2_else_and_439_nl;
  wire LOOPK2_else_and_441_nl;
  wire LOOPK2_else_and_443_nl;
  wire LOOPK2_else_and_445_nl;
  wire LOOPK2_else_and_447_nl;
  wire LOOPK2_else_and_449_nl;
  wire LOOPK2_else_and_451_nl;
  wire LOOPK2_else_and_453_nl;
  wire LOOPK2_else_and_455_nl;
  wire LOOPK2_else_and_457_nl;
  wire LOOPK2_else_and_459_nl;
  wire LOOPK2_else_and_461_nl;
  wire LOOPK2_else_and_463_nl;
  wire LOOPK2_else_and_465_nl;
  wire LOOPK2_else_and_467_nl;
  wire[37:0] LOOPK2_if_and_145_nl;
  wire LOOPK2_if_not_700_nl;
  wire LOOPK2_LOOPK2_nor_43_nl;
  wire LOOPK2_else_and_1513_nl;
  wire LOOPK2_else_and_1515_nl;
  wire LOOPK2_else_and_1517_nl;
  wire LOOPK2_else_and_1519_nl;
  wire LOOPK2_else_and_1521_nl;
  wire LOOPK2_else_and_1523_nl;
  wire LOOPK2_else_and_1525_nl;
  wire LOOPK2_else_and_1527_nl;
  wire LOOPK2_else_and_1529_nl;
  wire LOOPK2_else_and_1531_nl;
  wire LOOPK2_else_and_1533_nl;
  wire LOOPK2_else_and_1535_nl;
  wire LOOPK2_else_and_1537_nl;
  wire LOOPK2_else_and_1539_nl;
  wire LOOPK2_else_and_1541_nl;
  wire LOOPK2_else_and_1543_nl;
  wire LOOPK2_else_and_1545_nl;
  wire LOOPK2_else_and_1547_nl;
  wire[37:0] LOOPK2_if_and_144_nl;
  wire LOOPK2_if_not_718_nl;
  wire LOOPK2_LOOPK2_nor_14_nl;
  wire LOOPK2_else_and_469_nl;
  wire LOOPK2_else_and_471_nl;
  wire LOOPK2_else_and_473_nl;
  wire LOOPK2_else_and_475_nl;
  wire LOOPK2_else_and_477_nl;
  wire LOOPK2_else_and_479_nl;
  wire LOOPK2_else_and_481_nl;
  wire LOOPK2_else_and_483_nl;
  wire LOOPK2_else_and_485_nl;
  wire LOOPK2_else_and_487_nl;
  wire LOOPK2_else_and_489_nl;
  wire LOOPK2_else_and_491_nl;
  wire LOOPK2_else_and_493_nl;
  wire LOOPK2_else_and_495_nl;
  wire LOOPK2_else_and_497_nl;
  wire LOOPK2_else_and_499_nl;
  wire LOOPK2_else_and_501_nl;
  wire LOOPK2_else_and_503_nl;
  wire[37:0] LOOPK2_if_and_143_nl;
  wire LOOPK2_if_not_736_nl;
  wire LOOPK2_LOOPK2_nor_42_nl;
  wire LOOPK2_else_and_1477_nl;
  wire LOOPK2_else_and_1479_nl;
  wire LOOPK2_else_and_1481_nl;
  wire LOOPK2_else_and_1483_nl;
  wire LOOPK2_else_and_1485_nl;
  wire LOOPK2_else_and_1487_nl;
  wire LOOPK2_else_and_1489_nl;
  wire LOOPK2_else_and_1491_nl;
  wire LOOPK2_else_and_1493_nl;
  wire LOOPK2_else_and_1495_nl;
  wire LOOPK2_else_and_1497_nl;
  wire LOOPK2_else_and_1499_nl;
  wire LOOPK2_else_and_1501_nl;
  wire LOOPK2_else_and_1503_nl;
  wire LOOPK2_else_and_1505_nl;
  wire LOOPK2_else_and_1507_nl;
  wire LOOPK2_else_and_1509_nl;
  wire LOOPK2_else_and_1511_nl;
  wire[37:0] LOOPK2_if_and_142_nl;
  wire LOOPK2_if_not_754_nl;
  wire LOOPK2_LOOPK2_nor_15_nl;
  wire LOOPK2_else_and_505_nl;
  wire LOOPK2_else_and_507_nl;
  wire LOOPK2_else_and_509_nl;
  wire LOOPK2_else_and_511_nl;
  wire LOOPK2_else_and_513_nl;
  wire LOOPK2_else_and_515_nl;
  wire LOOPK2_else_and_517_nl;
  wire LOOPK2_else_and_519_nl;
  wire LOOPK2_else_and_521_nl;
  wire LOOPK2_else_and_523_nl;
  wire LOOPK2_else_and_525_nl;
  wire LOOPK2_else_and_527_nl;
  wire LOOPK2_else_and_529_nl;
  wire LOOPK2_else_and_531_nl;
  wire LOOPK2_else_and_533_nl;
  wire LOOPK2_else_and_535_nl;
  wire LOOPK2_else_and_537_nl;
  wire LOOPK2_else_and_539_nl;
  wire[37:0] LOOPK2_if_and_141_nl;
  wire LOOPK2_if_not_772_nl;
  wire LOOPK2_LOOPK2_nor_41_nl;
  wire LOOPK2_else_and_1441_nl;
  wire LOOPK2_else_and_1443_nl;
  wire LOOPK2_else_and_1445_nl;
  wire LOOPK2_else_and_1447_nl;
  wire LOOPK2_else_and_1449_nl;
  wire LOOPK2_else_and_1451_nl;
  wire LOOPK2_else_and_1453_nl;
  wire LOOPK2_else_and_1455_nl;
  wire LOOPK2_else_and_1457_nl;
  wire LOOPK2_else_and_1459_nl;
  wire LOOPK2_else_and_1461_nl;
  wire LOOPK2_else_and_1463_nl;
  wire LOOPK2_else_and_1465_nl;
  wire LOOPK2_else_and_1467_nl;
  wire LOOPK2_else_and_1469_nl;
  wire LOOPK2_else_and_1471_nl;
  wire LOOPK2_else_and_1473_nl;
  wire LOOPK2_else_and_1475_nl;
  wire[37:0] LOOPK2_if_and_140_nl;
  wire LOOPK2_if_not_790_nl;
  wire LOOPK2_LOOPK2_nor_16_nl;
  wire LOOPK2_else_and_541_nl;
  wire LOOPK2_else_and_543_nl;
  wire LOOPK2_else_and_545_nl;
  wire LOOPK2_else_and_547_nl;
  wire LOOPK2_else_and_549_nl;
  wire LOOPK2_else_and_551_nl;
  wire LOOPK2_else_and_553_nl;
  wire LOOPK2_else_and_555_nl;
  wire LOOPK2_else_and_557_nl;
  wire LOOPK2_else_and_559_nl;
  wire LOOPK2_else_and_561_nl;
  wire LOOPK2_else_and_563_nl;
  wire LOOPK2_else_and_565_nl;
  wire LOOPK2_else_and_567_nl;
  wire LOOPK2_else_and_569_nl;
  wire LOOPK2_else_and_571_nl;
  wire LOOPK2_else_and_573_nl;
  wire LOOPK2_else_and_575_nl;
  wire[37:0] LOOPK2_if_and_139_nl;
  wire LOOPK2_if_not_808_nl;
  wire LOOPK2_LOOPK2_nor_40_nl;
  wire LOOPK2_else_and_1405_nl;
  wire LOOPK2_else_and_1407_nl;
  wire LOOPK2_else_and_1409_nl;
  wire LOOPK2_else_and_1411_nl;
  wire LOOPK2_else_and_1413_nl;
  wire LOOPK2_else_and_1415_nl;
  wire LOOPK2_else_and_1417_nl;
  wire LOOPK2_else_and_1419_nl;
  wire LOOPK2_else_and_1421_nl;
  wire LOOPK2_else_and_1423_nl;
  wire LOOPK2_else_and_1425_nl;
  wire LOOPK2_else_and_1427_nl;
  wire LOOPK2_else_and_1429_nl;
  wire LOOPK2_else_and_1431_nl;
  wire LOOPK2_else_and_1433_nl;
  wire LOOPK2_else_and_1435_nl;
  wire LOOPK2_else_and_1437_nl;
  wire LOOPK2_else_and_1439_nl;
  wire[37:0] LOOPK2_if_and_138_nl;
  wire LOOPK2_if_not_826_nl;
  wire LOOPK2_LOOPK2_nor_17_nl;
  wire LOOPK2_else_and_577_nl;
  wire LOOPK2_else_and_579_nl;
  wire LOOPK2_else_and_581_nl;
  wire LOOPK2_else_and_583_nl;
  wire LOOPK2_else_and_585_nl;
  wire LOOPK2_else_and_587_nl;
  wire LOOPK2_else_and_589_nl;
  wire LOOPK2_else_and_591_nl;
  wire LOOPK2_else_and_593_nl;
  wire LOOPK2_else_and_595_nl;
  wire LOOPK2_else_and_597_nl;
  wire LOOPK2_else_and_599_nl;
  wire LOOPK2_else_and_601_nl;
  wire LOOPK2_else_and_603_nl;
  wire LOOPK2_else_and_605_nl;
  wire LOOPK2_else_and_607_nl;
  wire LOOPK2_else_and_609_nl;
  wire LOOPK2_else_and_611_nl;
  wire[37:0] LOOPK2_if_and_137_nl;
  wire LOOPK2_if_not_844_nl;
  wire LOOPK2_LOOPK2_nor_39_nl;
  wire LOOPK2_else_and_1369_nl;
  wire LOOPK2_else_and_1371_nl;
  wire LOOPK2_else_and_1373_nl;
  wire LOOPK2_else_and_1375_nl;
  wire LOOPK2_else_and_1377_nl;
  wire LOOPK2_else_and_1379_nl;
  wire LOOPK2_else_and_1381_nl;
  wire LOOPK2_else_and_1383_nl;
  wire LOOPK2_else_and_1385_nl;
  wire LOOPK2_else_and_1387_nl;
  wire LOOPK2_else_and_1389_nl;
  wire LOOPK2_else_and_1391_nl;
  wire LOOPK2_else_and_1393_nl;
  wire LOOPK2_else_and_1395_nl;
  wire LOOPK2_else_and_1397_nl;
  wire LOOPK2_else_and_1399_nl;
  wire LOOPK2_else_and_1401_nl;
  wire LOOPK2_else_and_1403_nl;
  wire[37:0] LOOPK2_if_and_136_nl;
  wire LOOPK2_if_not_862_nl;
  wire LOOPK2_LOOPK2_nor_18_nl;
  wire LOOPK2_else_and_613_nl;
  wire LOOPK2_else_and_615_nl;
  wire LOOPK2_else_and_617_nl;
  wire LOOPK2_else_and_619_nl;
  wire LOOPK2_else_and_621_nl;
  wire LOOPK2_else_and_623_nl;
  wire LOOPK2_else_and_625_nl;
  wire LOOPK2_else_and_627_nl;
  wire LOOPK2_else_and_629_nl;
  wire LOOPK2_else_and_631_nl;
  wire LOOPK2_else_and_633_nl;
  wire LOOPK2_else_and_635_nl;
  wire LOOPK2_else_and_637_nl;
  wire LOOPK2_else_and_639_nl;
  wire LOOPK2_else_and_641_nl;
  wire LOOPK2_else_and_643_nl;
  wire LOOPK2_else_and_645_nl;
  wire LOOPK2_else_and_647_nl;
  wire[37:0] LOOPK2_if_and_135_nl;
  wire LOOPK2_if_not_880_nl;
  wire LOOPK2_LOOPK2_nor_38_nl;
  wire LOOPK2_else_and_1333_nl;
  wire LOOPK2_else_and_1335_nl;
  wire LOOPK2_else_and_1337_nl;
  wire LOOPK2_else_and_1339_nl;
  wire LOOPK2_else_and_1341_nl;
  wire LOOPK2_else_and_1343_nl;
  wire LOOPK2_else_and_1345_nl;
  wire LOOPK2_else_and_1347_nl;
  wire LOOPK2_else_and_1349_nl;
  wire LOOPK2_else_and_1351_nl;
  wire LOOPK2_else_and_1353_nl;
  wire LOOPK2_else_and_1355_nl;
  wire LOOPK2_else_and_1357_nl;
  wire LOOPK2_else_and_1359_nl;
  wire LOOPK2_else_and_1361_nl;
  wire LOOPK2_else_and_1363_nl;
  wire LOOPK2_else_and_1365_nl;
  wire LOOPK2_else_and_1367_nl;
  wire[37:0] LOOPK2_if_and_134_nl;
  wire LOOPK2_if_not_898_nl;
  wire LOOPK2_LOOPK2_nor_19_nl;
  wire LOOPK2_else_and_649_nl;
  wire LOOPK2_else_and_651_nl;
  wire LOOPK2_else_and_653_nl;
  wire LOOPK2_else_and_655_nl;
  wire LOOPK2_else_and_657_nl;
  wire LOOPK2_else_and_659_nl;
  wire LOOPK2_else_and_661_nl;
  wire LOOPK2_else_and_663_nl;
  wire LOOPK2_else_and_665_nl;
  wire LOOPK2_else_and_667_nl;
  wire LOOPK2_else_and_669_nl;
  wire LOOPK2_else_and_671_nl;
  wire LOOPK2_else_and_673_nl;
  wire LOOPK2_else_and_675_nl;
  wire LOOPK2_else_and_677_nl;
  wire LOOPK2_else_and_679_nl;
  wire LOOPK2_else_and_681_nl;
  wire LOOPK2_else_and_683_nl;
  wire[37:0] LOOPK2_if_and_133_nl;
  wire LOOPK2_if_not_916_nl;
  wire LOOPK2_LOOPK2_nor_37_nl;
  wire LOOPK2_else_and_1297_nl;
  wire LOOPK2_else_and_1299_nl;
  wire LOOPK2_else_and_1301_nl;
  wire LOOPK2_else_and_1303_nl;
  wire LOOPK2_else_and_1305_nl;
  wire LOOPK2_else_and_1307_nl;
  wire LOOPK2_else_and_1309_nl;
  wire LOOPK2_else_and_1311_nl;
  wire LOOPK2_else_and_1313_nl;
  wire LOOPK2_else_and_1315_nl;
  wire LOOPK2_else_and_1317_nl;
  wire LOOPK2_else_and_1319_nl;
  wire LOOPK2_else_and_1321_nl;
  wire LOOPK2_else_and_1323_nl;
  wire LOOPK2_else_and_1325_nl;
  wire LOOPK2_else_and_1327_nl;
  wire LOOPK2_else_and_1329_nl;
  wire LOOPK2_else_and_1331_nl;
  wire[37:0] LOOPK2_if_and_132_nl;
  wire LOOPK2_if_not_934_nl;
  wire LOOPK2_LOOPK2_nor_20_nl;
  wire LOOPK2_else_and_685_nl;
  wire LOOPK2_else_and_687_nl;
  wire LOOPK2_else_and_689_nl;
  wire LOOPK2_else_and_691_nl;
  wire LOOPK2_else_and_693_nl;
  wire LOOPK2_else_and_695_nl;
  wire LOOPK2_else_and_697_nl;
  wire LOOPK2_else_and_699_nl;
  wire LOOPK2_else_and_701_nl;
  wire LOOPK2_else_and_703_nl;
  wire LOOPK2_else_and_705_nl;
  wire LOOPK2_else_and_707_nl;
  wire LOOPK2_else_and_709_nl;
  wire LOOPK2_else_and_711_nl;
  wire LOOPK2_else_and_713_nl;
  wire LOOPK2_else_and_715_nl;
  wire LOOPK2_else_and_717_nl;
  wire LOOPK2_else_and_719_nl;
  wire[37:0] LOOPK2_if_and_131_nl;
  wire LOOPK2_if_not_952_nl;
  wire LOOPK2_LOOPK2_nor_36_nl;
  wire LOOPK2_else_and_1261_nl;
  wire LOOPK2_else_and_1263_nl;
  wire LOOPK2_else_and_1265_nl;
  wire LOOPK2_else_and_1267_nl;
  wire LOOPK2_else_and_1269_nl;
  wire LOOPK2_else_and_1271_nl;
  wire LOOPK2_else_and_1273_nl;
  wire LOOPK2_else_and_1275_nl;
  wire LOOPK2_else_and_1277_nl;
  wire LOOPK2_else_and_1279_nl;
  wire LOOPK2_else_and_1281_nl;
  wire LOOPK2_else_and_1283_nl;
  wire LOOPK2_else_and_1285_nl;
  wire LOOPK2_else_and_1287_nl;
  wire LOOPK2_else_and_1289_nl;
  wire LOOPK2_else_and_1291_nl;
  wire LOOPK2_else_and_1293_nl;
  wire LOOPK2_else_and_1295_nl;
  wire[37:0] LOOPK2_if_and_130_nl;
  wire LOOPK2_if_not_970_nl;
  wire LOOPK2_LOOPK2_nor_21_nl;
  wire LOOPK2_else_and_721_nl;
  wire LOOPK2_else_and_723_nl;
  wire LOOPK2_else_and_725_nl;
  wire LOOPK2_else_and_727_nl;
  wire LOOPK2_else_and_729_nl;
  wire LOOPK2_else_and_731_nl;
  wire LOOPK2_else_and_733_nl;
  wire LOOPK2_else_and_735_nl;
  wire LOOPK2_else_and_737_nl;
  wire LOOPK2_else_and_739_nl;
  wire LOOPK2_else_and_741_nl;
  wire LOOPK2_else_and_743_nl;
  wire LOOPK2_else_and_745_nl;
  wire LOOPK2_else_and_747_nl;
  wire LOOPK2_else_and_749_nl;
  wire LOOPK2_else_and_751_nl;
  wire LOOPK2_else_and_753_nl;
  wire LOOPK2_else_and_755_nl;
  wire[37:0] LOOPK2_if_and_129_nl;
  wire LOOPK2_if_not_988_nl;
  wire LOOPK2_LOOPK2_nor_35_nl;
  wire LOOPK2_else_and_1225_nl;
  wire LOOPK2_else_and_1227_nl;
  wire LOOPK2_else_and_1229_nl;
  wire LOOPK2_else_and_1231_nl;
  wire LOOPK2_else_and_1233_nl;
  wire LOOPK2_else_and_1235_nl;
  wire LOOPK2_else_and_1237_nl;
  wire LOOPK2_else_and_1239_nl;
  wire LOOPK2_else_and_1241_nl;
  wire LOOPK2_else_and_1243_nl;
  wire LOOPK2_else_and_1245_nl;
  wire LOOPK2_else_and_1247_nl;
  wire LOOPK2_else_and_1249_nl;
  wire LOOPK2_else_and_1251_nl;
  wire LOOPK2_else_and_1253_nl;
  wire LOOPK2_else_and_1255_nl;
  wire LOOPK2_else_and_1257_nl;
  wire LOOPK2_else_and_1259_nl;
  wire[37:0] LOOPK2_if_and_128_nl;
  wire LOOPK2_if_not_1006_nl;
  wire LOOPK2_LOOPK2_nor_22_nl;
  wire LOOPK2_else_and_757_nl;
  wire LOOPK2_else_and_759_nl;
  wire LOOPK2_else_and_761_nl;
  wire LOOPK2_else_and_763_nl;
  wire LOOPK2_else_and_765_nl;
  wire LOOPK2_else_and_767_nl;
  wire LOOPK2_else_and_769_nl;
  wire LOOPK2_else_and_771_nl;
  wire LOOPK2_else_and_773_nl;
  wire LOOPK2_else_and_775_nl;
  wire LOOPK2_else_and_777_nl;
  wire LOOPK2_else_and_779_nl;
  wire LOOPK2_else_and_781_nl;
  wire LOOPK2_else_and_783_nl;
  wire LOOPK2_else_and_785_nl;
  wire LOOPK2_else_and_787_nl;
  wire LOOPK2_else_and_789_nl;
  wire LOOPK2_else_and_791_nl;
  wire[37:0] LOOPK2_if_and_127_nl;
  wire LOOPK2_if_not_1024_nl;
  wire LOOPK2_LOOPK2_nor_34_nl;
  wire LOOPK2_else_and_1189_nl;
  wire LOOPK2_else_and_1191_nl;
  wire LOOPK2_else_and_1193_nl;
  wire LOOPK2_else_and_1195_nl;
  wire LOOPK2_else_and_1197_nl;
  wire LOOPK2_else_and_1199_nl;
  wire LOOPK2_else_and_1201_nl;
  wire LOOPK2_else_and_1203_nl;
  wire LOOPK2_else_and_1205_nl;
  wire LOOPK2_else_and_1207_nl;
  wire LOOPK2_else_and_1209_nl;
  wire LOOPK2_else_and_1211_nl;
  wire LOOPK2_else_and_1213_nl;
  wire LOOPK2_else_and_1215_nl;
  wire LOOPK2_else_and_1217_nl;
  wire LOOPK2_else_and_1219_nl;
  wire LOOPK2_else_and_1221_nl;
  wire LOOPK2_else_and_1223_nl;
  wire[37:0] LOOPK2_if_and_126_nl;
  wire LOOPK2_if_not_1042_nl;
  wire LOOPK2_LOOPK2_nor_23_nl;
  wire LOOPK2_else_and_793_nl;
  wire LOOPK2_else_and_795_nl;
  wire LOOPK2_else_and_797_nl;
  wire LOOPK2_else_and_799_nl;
  wire LOOPK2_else_and_801_nl;
  wire LOOPK2_else_and_803_nl;
  wire LOOPK2_else_and_805_nl;
  wire LOOPK2_else_and_807_nl;
  wire LOOPK2_else_and_809_nl;
  wire LOOPK2_else_and_811_nl;
  wire LOOPK2_else_and_813_nl;
  wire LOOPK2_else_and_815_nl;
  wire LOOPK2_else_and_817_nl;
  wire LOOPK2_else_and_819_nl;
  wire LOOPK2_else_and_821_nl;
  wire LOOPK2_else_and_823_nl;
  wire LOOPK2_else_and_825_nl;
  wire LOOPK2_else_and_827_nl;
  wire[37:0] LOOPK2_if_and_125_nl;
  wire LOOPK2_if_not_1060_nl;
  wire LOOPK2_LOOPK2_nor_33_nl;
  wire LOOPK2_else_and_1153_nl;
  wire LOOPK2_else_and_1155_nl;
  wire LOOPK2_else_and_1157_nl;
  wire LOOPK2_else_and_1159_nl;
  wire LOOPK2_else_and_1161_nl;
  wire LOOPK2_else_and_1163_nl;
  wire LOOPK2_else_and_1165_nl;
  wire LOOPK2_else_and_1167_nl;
  wire LOOPK2_else_and_1169_nl;
  wire LOOPK2_else_and_1171_nl;
  wire LOOPK2_else_and_1173_nl;
  wire LOOPK2_else_and_1175_nl;
  wire LOOPK2_else_and_1177_nl;
  wire LOOPK2_else_and_1179_nl;
  wire LOOPK2_else_and_1181_nl;
  wire LOOPK2_else_and_1183_nl;
  wire LOOPK2_else_and_1185_nl;
  wire LOOPK2_else_and_1187_nl;
  wire[37:0] LOOPK2_if_and_124_nl;
  wire LOOPK2_if_not_1078_nl;
  wire LOOPK2_LOOPK2_nor_24_nl;
  wire LOOPK2_else_and_829_nl;
  wire LOOPK2_else_and_831_nl;
  wire LOOPK2_else_and_833_nl;
  wire LOOPK2_else_and_835_nl;
  wire LOOPK2_else_and_837_nl;
  wire LOOPK2_else_and_839_nl;
  wire LOOPK2_else_and_841_nl;
  wire LOOPK2_else_and_843_nl;
  wire LOOPK2_else_and_845_nl;
  wire LOOPK2_else_and_847_nl;
  wire LOOPK2_else_and_849_nl;
  wire LOOPK2_else_and_851_nl;
  wire LOOPK2_else_and_853_nl;
  wire LOOPK2_else_and_855_nl;
  wire LOOPK2_else_and_857_nl;
  wire LOOPK2_else_and_859_nl;
  wire LOOPK2_else_and_861_nl;
  wire LOOPK2_else_and_863_nl;
  wire[37:0] LOOPK2_if_and_123_nl;
  wire LOOPK2_if_not_1096_nl;
  wire LOOPK2_LOOPK2_nor_32_nl;
  wire LOOPK2_else_and_1117_nl;
  wire LOOPK2_else_and_1119_nl;
  wire LOOPK2_else_and_1121_nl;
  wire LOOPK2_else_and_1123_nl;
  wire LOOPK2_else_and_1125_nl;
  wire LOOPK2_else_and_1127_nl;
  wire LOOPK2_else_and_1129_nl;
  wire LOOPK2_else_and_1131_nl;
  wire LOOPK2_else_and_1133_nl;
  wire LOOPK2_else_and_1135_nl;
  wire LOOPK2_else_and_1137_nl;
  wire LOOPK2_else_and_1139_nl;
  wire LOOPK2_else_and_1141_nl;
  wire LOOPK2_else_and_1143_nl;
  wire LOOPK2_else_and_1145_nl;
  wire LOOPK2_else_and_1147_nl;
  wire LOOPK2_else_and_1149_nl;
  wire LOOPK2_else_and_1151_nl;
  wire[37:0] LOOPK2_if_and_122_nl;
  wire LOOPK2_if_not_1114_nl;
  wire LOOPK2_LOOPK2_nor_25_nl;
  wire LOOPK2_else_and_865_nl;
  wire LOOPK2_else_and_867_nl;
  wire LOOPK2_else_and_869_nl;
  wire LOOPK2_else_and_871_nl;
  wire LOOPK2_else_and_873_nl;
  wire LOOPK2_else_and_875_nl;
  wire LOOPK2_else_and_877_nl;
  wire LOOPK2_else_and_879_nl;
  wire LOOPK2_else_and_881_nl;
  wire LOOPK2_else_and_883_nl;
  wire LOOPK2_else_and_885_nl;
  wire LOOPK2_else_and_887_nl;
  wire LOOPK2_else_and_889_nl;
  wire LOOPK2_else_and_891_nl;
  wire LOOPK2_else_and_893_nl;
  wire LOOPK2_else_and_895_nl;
  wire LOOPK2_else_and_897_nl;
  wire LOOPK2_else_and_899_nl;
  wire[37:0] LOOPK2_if_and_121_nl;
  wire LOOPK2_if_not_1132_nl;
  wire LOOPK2_LOOPK2_nor_31_nl;
  wire LOOPK2_else_and_1081_nl;
  wire LOOPK2_else_and_1083_nl;
  wire LOOPK2_else_and_1085_nl;
  wire LOOPK2_else_and_1087_nl;
  wire LOOPK2_else_and_1089_nl;
  wire LOOPK2_else_and_1091_nl;
  wire LOOPK2_else_and_1093_nl;
  wire LOOPK2_else_and_1095_nl;
  wire LOOPK2_else_and_1097_nl;
  wire LOOPK2_else_and_1099_nl;
  wire LOOPK2_else_and_1101_nl;
  wire LOOPK2_else_and_1103_nl;
  wire LOOPK2_else_and_1105_nl;
  wire LOOPK2_else_and_1107_nl;
  wire LOOPK2_else_and_1109_nl;
  wire LOOPK2_else_and_1111_nl;
  wire LOOPK2_else_and_1113_nl;
  wire LOOPK2_else_and_1115_nl;
  wire[37:0] LOOPK2_if_and_120_nl;
  wire LOOPK2_if_not_1150_nl;
  wire LOOPK2_LOOPK2_nor_26_nl;
  wire LOOPK2_else_and_901_nl;
  wire LOOPK2_else_and_903_nl;
  wire LOOPK2_else_and_905_nl;
  wire LOOPK2_else_and_907_nl;
  wire LOOPK2_else_and_909_nl;
  wire LOOPK2_else_and_911_nl;
  wire LOOPK2_else_and_913_nl;
  wire LOOPK2_else_and_915_nl;
  wire LOOPK2_else_and_917_nl;
  wire LOOPK2_else_and_919_nl;
  wire LOOPK2_else_and_921_nl;
  wire LOOPK2_else_and_923_nl;
  wire LOOPK2_else_and_925_nl;
  wire LOOPK2_else_and_927_nl;
  wire LOOPK2_else_and_929_nl;
  wire LOOPK2_else_and_931_nl;
  wire LOOPK2_else_and_933_nl;
  wire LOOPK2_else_and_935_nl;
  wire[37:0] LOOPK2_if_and_119_nl;
  wire LOOPK2_if_not_1168_nl;
  wire LOOPK2_LOOPK2_nor_30_nl;
  wire LOOPK2_else_and_1045_nl;
  wire LOOPK2_else_and_1047_nl;
  wire LOOPK2_else_and_1049_nl;
  wire LOOPK2_else_and_1051_nl;
  wire LOOPK2_else_and_1053_nl;
  wire LOOPK2_else_and_1055_nl;
  wire LOOPK2_else_and_1057_nl;
  wire LOOPK2_else_and_1059_nl;
  wire LOOPK2_else_and_1061_nl;
  wire LOOPK2_else_and_1063_nl;
  wire LOOPK2_else_and_1065_nl;
  wire LOOPK2_else_and_1067_nl;
  wire LOOPK2_else_and_1069_nl;
  wire LOOPK2_else_and_1071_nl;
  wire LOOPK2_else_and_1073_nl;
  wire LOOPK2_else_and_1075_nl;
  wire LOOPK2_else_and_1077_nl;
  wire LOOPK2_else_and_1079_nl;
  wire[37:0] LOOPK2_if_and_118_nl;
  wire LOOPK2_if_not_1186_nl;
  wire LOOPK2_LOOPK2_nor_27_nl;
  wire LOOPK2_else_and_937_nl;
  wire LOOPK2_else_and_939_nl;
  wire LOOPK2_else_and_941_nl;
  wire LOOPK2_else_and_943_nl;
  wire LOOPK2_else_and_945_nl;
  wire LOOPK2_else_and_947_nl;
  wire LOOPK2_else_and_949_nl;
  wire LOOPK2_else_and_951_nl;
  wire LOOPK2_else_and_953_nl;
  wire LOOPK2_else_and_955_nl;
  wire LOOPK2_else_and_957_nl;
  wire LOOPK2_else_and_959_nl;
  wire LOOPK2_else_and_961_nl;
  wire LOOPK2_else_and_963_nl;
  wire LOOPK2_else_and_965_nl;
  wire LOOPK2_else_and_967_nl;
  wire LOOPK2_else_and_969_nl;
  wire LOOPK2_else_and_971_nl;
  wire[37:0] LOOPK2_if_and_117_nl;
  wire LOOPK2_if_not_1204_nl;
  wire LOOPK2_LOOPK2_nor_29_nl;
  wire LOOPK2_else_and_1009_nl;
  wire LOOPK2_else_and_1011_nl;
  wire LOOPK2_else_and_1013_nl;
  wire LOOPK2_else_and_1015_nl;
  wire LOOPK2_else_and_1017_nl;
  wire LOOPK2_else_and_1019_nl;
  wire LOOPK2_else_and_1021_nl;
  wire LOOPK2_else_and_1023_nl;
  wire LOOPK2_else_and_1025_nl;
  wire LOOPK2_else_and_1027_nl;
  wire LOOPK2_else_and_1029_nl;
  wire LOOPK2_else_and_1031_nl;
  wire LOOPK2_else_and_1033_nl;
  wire LOOPK2_else_and_1035_nl;
  wire LOOPK2_else_and_1037_nl;
  wire LOOPK2_else_and_1039_nl;
  wire LOOPK2_else_and_1041_nl;
  wire LOOPK2_else_and_1043_nl;
  wire[37:0] LOOPK2_if_and_116_nl;
  wire LOOPK2_if_not_1222_nl;
  wire LOOPK2_LOOPK2_nor_28_nl;
  wire LOOPK2_else_and_973_nl;
  wire LOOPK2_else_and_975_nl;
  wire LOOPK2_else_and_977_nl;
  wire LOOPK2_else_and_979_nl;
  wire LOOPK2_else_and_981_nl;
  wire LOOPK2_else_and_983_nl;
  wire LOOPK2_else_and_985_nl;
  wire LOOPK2_else_and_987_nl;
  wire LOOPK2_else_and_989_nl;
  wire LOOPK2_else_and_991_nl;
  wire LOOPK2_else_and_993_nl;
  wire LOOPK2_else_and_995_nl;
  wire LOOPK2_else_and_997_nl;
  wire LOOPK2_else_and_999_nl;
  wire LOOPK2_else_and_1001_nl;
  wire LOOPK2_else_and_1003_nl;
  wire LOOPK2_else_and_1005_nl;
  wire LOOPK2_else_and_1007_nl;
  wire[36:0] operator_38_true_acc_nl;
  wire[37:0] nl_operator_38_true_acc_nl;
  wire[35:0] operator_38_true_operator_38_true_mux_nl;
  wire or_1731_nl;
  wire[5:0] operator_6_false_3_mux_1_nl;
  wire or_1746_nl;
  wire operator_8_false_operator_8_false_and_1_nl;
  wire operator_8_false_mux_3_nl;
  wire[5:0] operator_8_false_mux_4_nl;
  wire operator_8_false_operator_8_false_or_1_nl;
  wire operator_7_false_1_operator_7_false_1_and_1_nl;
  wire[5:0] operator_7_false_1_mux_2_nl;
  wire[15:0] LOOPK2_mux_172_nl;
  wire[15:0] LOOPK2_mux_173_nl;
  wire[15:0] LOOPK2_LOOPK2_mux_1_nl;
  wire LOOPL1_LOOPL1_and_2_nl;
  wire LOOPL1_mux_66_nl;
  wire[15:0] LOOPL1_mux1h_4_nl;
  wire[37:0] LOOPL1_mux1h_5_nl;
  wire[31:0] LOOPL2_LOOPL2_mux_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr0;
  assign nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr0 = LOOPL1_LOOPL1_and_tmp
      & nor_169_cse;
  wire  nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr1;
  assign nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr1 = ~
      nor_169_cse;
  wire mux_5_nl;
  wire  nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPK3_C_0_tr0;
  assign mux_5_nl = MUX_s_1_2_2((~ LOOPK3_if_unequal_tmp), LOOPK3_if_equal_tmp, z_out_2[0]);
  assign nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPK3_C_0_tr0 = mux_5_nl
      & (~ (z_out_2[7]));
  wire  nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL2_C_0_tr0;
  assign nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL2_C_0_tr0 = LOOPL2_l_sva
      == conv_s2s_8_32(z_out_2);
  ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci ATTENTION_IP_Attention_Calculator_run_q_chan2_rsci_inst
      (
      .q_chan2_rsc_dat(q_chan2_rsc_dat),
      .q_chan2_rsc_vld(q_chan2_rsc_vld),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy),
      .q_chan2_rsci_oswt(reg_q_chan2_rsci_oswt_cse),
      .q_chan2_rsci_wen_comp(q_chan2_rsci_wen_comp),
      .q_chan2_rsci_idat_mxwt(q_chan2_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci ATTENTION_IP_Attention_Calculator_run_k_chan2_rsci_inst
      (
      .k_chan2_rsc_dat(k_chan2_rsc_dat),
      .k_chan2_rsc_vld(k_chan2_rsc_vld),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy),
      .k_chan2_rsci_oswt(reg_k_chan2_rsci_oswt_cse),
      .k_chan2_rsci_wen_comp(k_chan2_rsci_wen_comp),
      .k_chan2_rsci_idat_mxwt(k_chan2_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci ATTENTION_IP_Attention_Calculator_run_v_chan2_rsci_inst
      (
      .v_chan2_rsc_dat(v_chan2_rsc_dat),
      .v_chan2_rsc_vld(v_chan2_rsc_vld),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy),
      .v_chan2_rsci_oswt(reg_v_chan2_rsci_oswt_cse),
      .v_chan2_rsci_wen_comp(v_chan2_rsci_wen_comp),
      .v_chan2_rsci_idat_mxwt(v_chan2_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci ATTENTION_IP_Attention_Calculator_run_dout_chan_rsci_inst
      (
      .dout_chan_rsc_dat(dout_chan_rsc_dat),
      .dout_chan_rsc_vld(dout_chan_rsc_vld),
      .dout_chan_rsc_rdy(dout_chan_rsc_rdy),
      .dout_chan_rsci_oswt(reg_dout_chan_rsci_oswt_cse),
      .dout_chan_rsci_wen_comp(dout_chan_rsci_wen_comp),
      .dout_chan_rsci_idat(dout_chan_rsci_idat)
    );
  ATTENTION_IP_Attention_Calculator_run_staller ATTENTION_IP_Attention_Calculator_run_staller_inst
      (
      .run_wen(run_wen),
      .q_chan2_rsci_wen_comp(q_chan2_rsci_wen_comp),
      .k_chan2_rsci_wen_comp(k_chan2_rsci_wen_comp),
      .v_chan2_rsci_wen_comp(v_chan2_rsci_wen_comp),
      .dout_chan_rsci_wen_comp(dout_chan_rsci_wen_comp)
    );
  ATTENTION_IP_Attention_Calculator_run_run_fsm ATTENTION_IP_Attention_Calculator_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .LOOPL1_C_0_tr0(nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr0),
      .LOOPL1_C_0_tr1(nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL1_C_0_tr1),
      .LOOPK2_C_0_tr0(LOOPK4_LOOPK4_if_1_and_tmp),
      .LOOPK3_C_0_tr0(nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPK3_C_0_tr0),
      .LOOPL2_C_0_tr0(nl_ATTENTION_IP_Attention_Calculator_run_run_fsm_inst_LOOPL2_C_0_tr0),
      .LOOPK4_C_1_tr0(LOOPK4_LOOPK4_if_1_and_tmp),
      .LOOPK5_C_1_tr0(LOOPK1_endflag_sva),
      .LOOPJ1_C_3_tr0(LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp),
      .LOOPI1_C_0_tr0(LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp)
    );
  assign LOOPI1_i_or_cse = (fsm_output[0]) | (fsm_output[15]);
  assign nand_22_cse = ~((fsm_output[7]) & (LOOPK5_k_sva_5_0[4:0]==5'b01111));
  assign nand_31_cse = ~((fsm_output[7]) & (LOOPK5_k_sva_5_0[3:0]==4'b0111));
  assign nand_34_cse = ~((LOOPK5_k_sva_5_0[4:3]==2'b11));
  assign nand_44_cse = ~((fsm_output[7]) & (LOOPK5_k_sva_5_0[2:0]==3'b011));
  assign nand_47_cse = ~((LOOPK5_k_sva_5_0[4:2]==3'b111));
  assign nand_55_cse = ~((LOOPL2_l_sva[5:2]==4'b1111) & (fsm_output[10]));
  assign nand_58_cse = ~((LOOPL2_l_sva[5]) & (fsm_output[10]));
  assign nand_75_cse = ~((LOOPL2_l_sva[5:4]==2'b11) & (fsm_output[10]));
  assign nand_84_cse = ~((LOOPL2_l_sva[5:3]==3'b111) & (fsm_output[10]));
  assign or_1735_cse = (z_out_2[0]) | (z_out_2[7]) | LOOPK3_if_unequal_tmp;
  assign nor_14_cse = ~(LOOPK3_if_unequal_tmp | (z_out_2[7]) | (z_out_2[0]));
  assign and_2155_cse = (fsm_output[8]) & LOOPK1_endflag_sva;
  assign nor_169_cse = ~(LOOPL1_if_1_unequal_1_itm | (z_out_2[7]));
  assign nl_LOOPK1_acc_1_nl = conv_s2u_38_39(maxn_sva) - conv_s2u_13_39(LOOPL1_ac_int_cctor_sva[37:25]);
  assign LOOPK1_acc_1_nl = nl_LOOPK1_acc_1_nl[38:0];
  assign and_1639_rgt = (readslicef_39_1_38(LOOPK1_acc_1_nl)) & (fsm_output[4]);
  assign and_2169_cse = (~((fsm_output[8]) | (fsm_output[6]))) & (~((fsm_output[7])
      | (fsm_output[3])));
  assign nor_178_cse = ~((LOOPK5_k_sva_5_0[5:4]!=2'b00));
  assign nor_177_cse = ~((LOOPK5_k_sva_5_0[0]) | (LOOPK5_k_sva_5_0[2]) | (LOOPK5_k_sva_5_0[3]));
  assign nor_174_cse = ~((~ and_2169_cse) | (LOOPK5_k_sva_5_0[1]));
  assign nor_240_cse = ~((LOOPK5_k_sva_5_0[0]) | (LOOPK5_k_sva_5_0[2]));
  assign LOOPK5_k_nor_seb = ~((fsm_output[16]) | (fsm_output[2]) | (fsm_output[14])
      | (fsm_output[1]) | LOOPI1_i_or_cse | (fsm_output[4]) | (LOOPK4_LOOPK4_if_1_and_tmp
      & (fsm_output[11])));
  assign LOOPK1_and_61_cse = run_wen & (~(LOOPK1_endflag_sva & LOOPL1_LOOPL1_nor_tmp))
      & nor_169_cse;
  assign LOOPK2_if_not_232_nl = ~ LOOPK2_and_115_cse_sva_1;
  assign LOOPK2_if_and_171_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_55_lpi_5, LOOPK2_if_not_232_nl);
  assign LOOPK2_LOOPK2_nor_56_nl = ~((~(((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_115_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_115_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1981_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1983_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1985_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1987_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1989_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1991_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1993_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1995_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1997_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1999_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2001_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2003_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2005_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2007_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2009_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2011_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2013_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_2015_nl = LOOPK2_and_115_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_55_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_55_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_171_nl, {LOOPK2_LOOPK2_nor_56_nl , LOOPK2_else_and_1981_nl ,
      LOOPK2_else_and_1983_nl , LOOPK2_else_and_1985_nl , LOOPK2_else_and_1987_nl
      , LOOPK2_else_and_1989_nl , LOOPK2_else_and_1991_nl , LOOPK2_else_and_1993_nl
      , LOOPK2_else_and_1995_nl , LOOPK2_else_and_1997_nl , LOOPK2_else_and_1999_nl
      , LOOPK2_else_and_2001_nl , LOOPK2_else_and_2003_nl , LOOPK2_else_and_2005_nl
      , LOOPK2_else_and_2007_nl , LOOPK2_else_and_2009_nl , LOOPK2_else_and_2011_nl
      , LOOPK2_else_and_2013_nl , LOOPK2_else_and_2015_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_250_nl = ~ LOOPK2_and_114_cse_sva_1;
  assign LOOPK2_if_and_170_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_0_lpi_5, LOOPK2_if_not_250_nl);
  assign LOOPK2_LOOPK2_nor_1_nl = ~((~(((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_114_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_114_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_or_tmp_3 &
      (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_3_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_or_tmp_2 &
      (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_5_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_7_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_9_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_11_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_13_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_15_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_17_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_19_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_21_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_23_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_25_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_27_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_29_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_31_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_33_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_35_nl = LOOPK2_and_114_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_0_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_0_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_170_nl, {LOOPK2_LOOPK2_nor_1_nl , LOOPK2_else_and_1_nl , LOOPK2_else_and_3_nl
      , LOOPK2_else_and_5_nl , LOOPK2_else_and_7_nl , LOOPK2_else_and_9_nl , LOOPK2_else_and_11_nl
      , LOOPK2_else_and_13_nl , LOOPK2_else_and_15_nl , LOOPK2_else_and_17_nl , LOOPK2_else_and_19_nl
      , LOOPK2_else_and_21_nl , LOOPK2_else_and_23_nl , LOOPK2_else_and_25_nl , LOOPK2_else_and_27_nl
      , LOOPK2_else_and_29_nl , LOOPK2_else_and_31_nl , LOOPK2_else_and_33_nl , LOOPK2_else_and_35_nl
      , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_268_nl = ~ LOOPK2_and_113_cse_sva_1;
  assign LOOPK2_if_and_169_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_54_lpi_5, LOOPK2_if_not_268_nl);
  assign LOOPK2_LOOPK2_nor_55_nl = ~((~(((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_113_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_113_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1945_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1947_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1949_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1951_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1953_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1955_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1957_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1959_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1961_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1963_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1965_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1967_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1969_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1971_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1973_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1975_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1977_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1979_nl = LOOPK2_and_113_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_54_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_54_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_169_nl, {LOOPK2_LOOPK2_nor_55_nl , LOOPK2_else_and_1945_nl ,
      LOOPK2_else_and_1947_nl , LOOPK2_else_and_1949_nl , LOOPK2_else_and_1951_nl
      , LOOPK2_else_and_1953_nl , LOOPK2_else_and_1955_nl , LOOPK2_else_and_1957_nl
      , LOOPK2_else_and_1959_nl , LOOPK2_else_and_1961_nl , LOOPK2_else_and_1963_nl
      , LOOPK2_else_and_1965_nl , LOOPK2_else_and_1967_nl , LOOPK2_else_and_1969_nl
      , LOOPK2_else_and_1971_nl , LOOPK2_else_and_1973_nl , LOOPK2_else_and_1975_nl
      , LOOPK2_else_and_1977_nl , LOOPK2_else_and_1979_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_286_nl = ~ LOOPK2_and_112_cse_sva_1;
  assign LOOPK2_if_and_168_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_1_lpi_5, LOOPK2_if_not_286_nl);
  assign LOOPK2_LOOPK2_nor_2_nl = ~((~(((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_112_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_112_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_37_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_39_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_41_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_43_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_45_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_47_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_49_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_51_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_53_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_55_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_57_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_59_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_61_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_63_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_65_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_67_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_69_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_71_nl = LOOPK2_and_112_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_1_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_1_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_168_nl, {LOOPK2_LOOPK2_nor_2_nl , LOOPK2_else_and_37_nl , LOOPK2_else_and_39_nl
      , LOOPK2_else_and_41_nl , LOOPK2_else_and_43_nl , LOOPK2_else_and_45_nl , LOOPK2_else_and_47_nl
      , LOOPK2_else_and_49_nl , LOOPK2_else_and_51_nl , LOOPK2_else_and_53_nl , LOOPK2_else_and_55_nl
      , LOOPK2_else_and_57_nl , LOOPK2_else_and_59_nl , LOOPK2_else_and_61_nl , LOOPK2_else_and_63_nl
      , LOOPK2_else_and_65_nl , LOOPK2_else_and_67_nl , LOOPK2_else_and_69_nl , LOOPK2_else_and_71_nl
      , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_304_nl = ~ LOOPK2_and_111_cse_sva_1;
  assign LOOPK2_if_and_167_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_53_lpi_5, LOOPK2_if_not_304_nl);
  assign LOOPK2_LOOPK2_nor_54_nl = ~((~(((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_111_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_111_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1909_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1911_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1913_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1915_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1917_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1919_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1921_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1923_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1925_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1927_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1929_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1931_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1933_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1935_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1937_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1939_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1941_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1943_nl = LOOPK2_and_111_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_53_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_53_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_167_nl, {LOOPK2_LOOPK2_nor_54_nl , LOOPK2_else_and_1909_nl ,
      LOOPK2_else_and_1911_nl , LOOPK2_else_and_1913_nl , LOOPK2_else_and_1915_nl
      , LOOPK2_else_and_1917_nl , LOOPK2_else_and_1919_nl , LOOPK2_else_and_1921_nl
      , LOOPK2_else_and_1923_nl , LOOPK2_else_and_1925_nl , LOOPK2_else_and_1927_nl
      , LOOPK2_else_and_1929_nl , LOOPK2_else_and_1931_nl , LOOPK2_else_and_1933_nl
      , LOOPK2_else_and_1935_nl , LOOPK2_else_and_1937_nl , LOOPK2_else_and_1939_nl
      , LOOPK2_else_and_1941_nl , LOOPK2_else_and_1943_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_322_nl = ~ LOOPK2_and_110_cse_sva_1;
  assign LOOPK2_if_and_166_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_2_lpi_5, LOOPK2_if_not_322_nl);
  assign LOOPK2_LOOPK2_nor_3_nl = ~((~(((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_110_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_110_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_73_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_75_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_77_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_79_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_81_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_83_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_85_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_87_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_89_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_91_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_93_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_95_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_97_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_99_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_101_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_103_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_105_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_107_nl = LOOPK2_and_110_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_2_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_2_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_166_nl, {LOOPK2_LOOPK2_nor_3_nl , LOOPK2_else_and_73_nl , LOOPK2_else_and_75_nl
      , LOOPK2_else_and_77_nl , LOOPK2_else_and_79_nl , LOOPK2_else_and_81_nl , LOOPK2_else_and_83_nl
      , LOOPK2_else_and_85_nl , LOOPK2_else_and_87_nl , LOOPK2_else_and_89_nl , LOOPK2_else_and_91_nl
      , LOOPK2_else_and_93_nl , LOOPK2_else_and_95_nl , LOOPK2_else_and_97_nl , LOOPK2_else_and_99_nl
      , LOOPK2_else_and_101_nl , LOOPK2_else_and_103_nl , LOOPK2_else_and_105_nl
      , LOOPK2_else_and_107_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_340_nl = ~ LOOPK2_and_109_cse_sva_1;
  assign LOOPK2_if_and_165_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_52_lpi_5, LOOPK2_if_not_340_nl);
  assign LOOPK2_LOOPK2_nor_53_nl = ~((~(((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_109_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_109_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1873_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1875_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1877_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1879_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1881_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1883_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1885_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1887_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1889_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1891_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1893_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1895_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1897_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1899_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1901_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1903_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1905_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1907_nl = LOOPK2_and_109_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_52_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_52_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_165_nl, {LOOPK2_LOOPK2_nor_53_nl , LOOPK2_else_and_1873_nl ,
      LOOPK2_else_and_1875_nl , LOOPK2_else_and_1877_nl , LOOPK2_else_and_1879_nl
      , LOOPK2_else_and_1881_nl , LOOPK2_else_and_1883_nl , LOOPK2_else_and_1885_nl
      , LOOPK2_else_and_1887_nl , LOOPK2_else_and_1889_nl , LOOPK2_else_and_1891_nl
      , LOOPK2_else_and_1893_nl , LOOPK2_else_and_1895_nl , LOOPK2_else_and_1897_nl
      , LOOPK2_else_and_1899_nl , LOOPK2_else_and_1901_nl , LOOPK2_else_and_1903_nl
      , LOOPK2_else_and_1905_nl , LOOPK2_else_and_1907_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_358_nl = ~ LOOPK2_and_108_cse_sva_1;
  assign LOOPK2_if_and_164_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_3_lpi_5, LOOPK2_if_not_358_nl);
  assign LOOPK2_LOOPK2_nor_4_nl = ~((~(((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_108_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_108_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_109_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_111_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_113_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_115_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_117_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_119_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_121_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_123_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_125_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_127_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_129_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_131_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_133_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_135_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_137_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_139_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_141_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_143_nl = LOOPK2_and_108_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_3_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_3_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_164_nl, {LOOPK2_LOOPK2_nor_4_nl , LOOPK2_else_and_109_nl , LOOPK2_else_and_111_nl
      , LOOPK2_else_and_113_nl , LOOPK2_else_and_115_nl , LOOPK2_else_and_117_nl
      , LOOPK2_else_and_119_nl , LOOPK2_else_and_121_nl , LOOPK2_else_and_123_nl
      , LOOPK2_else_and_125_nl , LOOPK2_else_and_127_nl , LOOPK2_else_and_129_nl
      , LOOPK2_else_and_131_nl , LOOPK2_else_and_133_nl , LOOPK2_else_and_135_nl
      , LOOPK2_else_and_137_nl , LOOPK2_else_and_139_nl , LOOPK2_else_and_141_nl
      , LOOPK2_else_and_143_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_376_nl = ~ LOOPK2_and_107_cse_sva_1;
  assign LOOPK2_if_and_163_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_51_lpi_5, LOOPK2_if_not_376_nl);
  assign LOOPK2_LOOPK2_nor_52_nl = ~((~(((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_107_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_107_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1837_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1839_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1841_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1843_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1845_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1847_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1849_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1851_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1853_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1855_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1857_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1859_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1861_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1863_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1865_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1867_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1869_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1871_nl = LOOPK2_and_107_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_51_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_51_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_163_nl, {LOOPK2_LOOPK2_nor_52_nl , LOOPK2_else_and_1837_nl ,
      LOOPK2_else_and_1839_nl , LOOPK2_else_and_1841_nl , LOOPK2_else_and_1843_nl
      , LOOPK2_else_and_1845_nl , LOOPK2_else_and_1847_nl , LOOPK2_else_and_1849_nl
      , LOOPK2_else_and_1851_nl , LOOPK2_else_and_1853_nl , LOOPK2_else_and_1855_nl
      , LOOPK2_else_and_1857_nl , LOOPK2_else_and_1859_nl , LOOPK2_else_and_1861_nl
      , LOOPK2_else_and_1863_nl , LOOPK2_else_and_1865_nl , LOOPK2_else_and_1867_nl
      , LOOPK2_else_and_1869_nl , LOOPK2_else_and_1871_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_394_nl = ~ LOOPK2_and_106_cse_sva_1;
  assign LOOPK2_if_and_162_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_4_lpi_5, LOOPK2_if_not_394_nl);
  assign LOOPK2_LOOPK2_nor_5_nl = ~((~(((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_106_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_106_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_145_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_147_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_149_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_151_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_153_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_155_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_157_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_159_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_161_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_163_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_165_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_167_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_169_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_171_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_173_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_175_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_177_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_179_nl = LOOPK2_and_106_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_4_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_4_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_162_nl, {LOOPK2_LOOPK2_nor_5_nl , LOOPK2_else_and_145_nl , LOOPK2_else_and_147_nl
      , LOOPK2_else_and_149_nl , LOOPK2_else_and_151_nl , LOOPK2_else_and_153_nl
      , LOOPK2_else_and_155_nl , LOOPK2_else_and_157_nl , LOOPK2_else_and_159_nl
      , LOOPK2_else_and_161_nl , LOOPK2_else_and_163_nl , LOOPK2_else_and_165_nl
      , LOOPK2_else_and_167_nl , LOOPK2_else_and_169_nl , LOOPK2_else_and_171_nl
      , LOOPK2_else_and_173_nl , LOOPK2_else_and_175_nl , LOOPK2_else_and_177_nl
      , LOOPK2_else_and_179_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_412_nl = ~ LOOPK2_and_105_cse_sva_1;
  assign LOOPK2_if_and_161_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_50_lpi_5, LOOPK2_if_not_412_nl);
  assign LOOPK2_LOOPK2_nor_51_nl = ~((~(((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_105_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_105_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1801_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1803_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1805_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1807_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1809_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1811_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1813_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1815_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1817_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1819_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1821_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1823_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1825_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1827_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1829_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1831_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1833_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1835_nl = LOOPK2_and_105_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_50_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_50_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_161_nl, {LOOPK2_LOOPK2_nor_51_nl , LOOPK2_else_and_1801_nl ,
      LOOPK2_else_and_1803_nl , LOOPK2_else_and_1805_nl , LOOPK2_else_and_1807_nl
      , LOOPK2_else_and_1809_nl , LOOPK2_else_and_1811_nl , LOOPK2_else_and_1813_nl
      , LOOPK2_else_and_1815_nl , LOOPK2_else_and_1817_nl , LOOPK2_else_and_1819_nl
      , LOOPK2_else_and_1821_nl , LOOPK2_else_and_1823_nl , LOOPK2_else_and_1825_nl
      , LOOPK2_else_and_1827_nl , LOOPK2_else_and_1829_nl , LOOPK2_else_and_1831_nl
      , LOOPK2_else_and_1833_nl , LOOPK2_else_and_1835_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_430_nl = ~ LOOPK2_and_104_cse_sva_1;
  assign LOOPK2_if_and_160_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_5_lpi_5, LOOPK2_if_not_430_nl);
  assign LOOPK2_LOOPK2_nor_6_nl = ~((~(((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_104_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_104_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_181_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_183_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_185_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_187_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_189_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_191_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_193_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_195_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_197_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_199_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_201_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_203_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_205_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_207_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_209_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_211_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_213_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_215_nl = LOOPK2_and_104_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_5_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_5_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_160_nl, {LOOPK2_LOOPK2_nor_6_nl , LOOPK2_else_and_181_nl , LOOPK2_else_and_183_nl
      , LOOPK2_else_and_185_nl , LOOPK2_else_and_187_nl , LOOPK2_else_and_189_nl
      , LOOPK2_else_and_191_nl , LOOPK2_else_and_193_nl , LOOPK2_else_and_195_nl
      , LOOPK2_else_and_197_nl , LOOPK2_else_and_199_nl , LOOPK2_else_and_201_nl
      , LOOPK2_else_and_203_nl , LOOPK2_else_and_205_nl , LOOPK2_else_and_207_nl
      , LOOPK2_else_and_209_nl , LOOPK2_else_and_211_nl , LOOPK2_else_and_213_nl
      , LOOPK2_else_and_215_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_448_nl = ~ LOOPK2_and_103_cse_sva_1;
  assign LOOPK2_if_and_159_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_49_lpi_5, LOOPK2_if_not_448_nl);
  assign LOOPK2_LOOPK2_nor_50_nl = ~((~(((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_103_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_103_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1765_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1767_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1769_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1771_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1773_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1775_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1777_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1779_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1781_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1783_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1785_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1787_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1789_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1791_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1793_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1795_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1797_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1799_nl = LOOPK2_and_103_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_49_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_49_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_159_nl, {LOOPK2_LOOPK2_nor_50_nl , LOOPK2_else_and_1765_nl ,
      LOOPK2_else_and_1767_nl , LOOPK2_else_and_1769_nl , LOOPK2_else_and_1771_nl
      , LOOPK2_else_and_1773_nl , LOOPK2_else_and_1775_nl , LOOPK2_else_and_1777_nl
      , LOOPK2_else_and_1779_nl , LOOPK2_else_and_1781_nl , LOOPK2_else_and_1783_nl
      , LOOPK2_else_and_1785_nl , LOOPK2_else_and_1787_nl , LOOPK2_else_and_1789_nl
      , LOOPK2_else_and_1791_nl , LOOPK2_else_and_1793_nl , LOOPK2_else_and_1795_nl
      , LOOPK2_else_and_1797_nl , LOOPK2_else_and_1799_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_466_nl = ~ LOOPK2_and_102_cse_sva_1;
  assign LOOPK2_if_and_158_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_6_lpi_5, LOOPK2_if_not_466_nl);
  assign LOOPK2_LOOPK2_nor_7_nl = ~((~(((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_102_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_102_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_217_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_219_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_221_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_223_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_225_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_227_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_229_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_231_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_233_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_235_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_237_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_239_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_241_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_243_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_245_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_247_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_249_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_251_nl = LOOPK2_and_102_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_6_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_6_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_158_nl, {LOOPK2_LOOPK2_nor_7_nl , LOOPK2_else_and_217_nl , LOOPK2_else_and_219_nl
      , LOOPK2_else_and_221_nl , LOOPK2_else_and_223_nl , LOOPK2_else_and_225_nl
      , LOOPK2_else_and_227_nl , LOOPK2_else_and_229_nl , LOOPK2_else_and_231_nl
      , LOOPK2_else_and_233_nl , LOOPK2_else_and_235_nl , LOOPK2_else_and_237_nl
      , LOOPK2_else_and_239_nl , LOOPK2_else_and_241_nl , LOOPK2_else_and_243_nl
      , LOOPK2_else_and_245_nl , LOOPK2_else_and_247_nl , LOOPK2_else_and_249_nl
      , LOOPK2_else_and_251_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_484_nl = ~ LOOPK2_and_101_cse_sva_1;
  assign LOOPK2_if_and_157_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_48_lpi_5, LOOPK2_if_not_484_nl);
  assign LOOPK2_LOOPK2_nor_49_nl = ~((~(((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_101_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_101_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1729_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1731_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1733_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1735_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1737_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1739_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1741_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1743_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1745_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1747_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1749_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1751_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1753_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1755_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1757_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1759_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1761_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1763_nl = LOOPK2_and_101_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_48_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_48_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_157_nl, {LOOPK2_LOOPK2_nor_49_nl , LOOPK2_else_and_1729_nl ,
      LOOPK2_else_and_1731_nl , LOOPK2_else_and_1733_nl , LOOPK2_else_and_1735_nl
      , LOOPK2_else_and_1737_nl , LOOPK2_else_and_1739_nl , LOOPK2_else_and_1741_nl
      , LOOPK2_else_and_1743_nl , LOOPK2_else_and_1745_nl , LOOPK2_else_and_1747_nl
      , LOOPK2_else_and_1749_nl , LOOPK2_else_and_1751_nl , LOOPK2_else_and_1753_nl
      , LOOPK2_else_and_1755_nl , LOOPK2_else_and_1757_nl , LOOPK2_else_and_1759_nl
      , LOOPK2_else_and_1761_nl , LOOPK2_else_and_1763_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_502_nl = ~ LOOPK2_and_100_cse_sva_1;
  assign LOOPK2_if_and_156_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_7_lpi_5, LOOPK2_if_not_502_nl);
  assign LOOPK2_LOOPK2_nor_8_nl = ~((~(((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_100_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_100_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_253_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_255_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_257_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_259_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_261_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_263_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_265_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_267_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_269_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_271_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_273_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_275_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_277_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_279_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_281_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_283_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_285_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_287_nl = LOOPK2_and_100_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_7_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_7_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_156_nl, {LOOPK2_LOOPK2_nor_8_nl , LOOPK2_else_and_253_nl , LOOPK2_else_and_255_nl
      , LOOPK2_else_and_257_nl , LOOPK2_else_and_259_nl , LOOPK2_else_and_261_nl
      , LOOPK2_else_and_263_nl , LOOPK2_else_and_265_nl , LOOPK2_else_and_267_nl
      , LOOPK2_else_and_269_nl , LOOPK2_else_and_271_nl , LOOPK2_else_and_273_nl
      , LOOPK2_else_and_275_nl , LOOPK2_else_and_277_nl , LOOPK2_else_and_279_nl
      , LOOPK2_else_and_281_nl , LOOPK2_else_and_283_nl , LOOPK2_else_and_285_nl
      , LOOPK2_else_and_287_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_520_nl = ~ LOOPK2_and_99_cse_sva_1;
  assign LOOPK2_if_and_155_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_47_lpi_5, LOOPK2_if_not_520_nl);
  assign LOOPK2_LOOPK2_nor_48_nl = ~((~(((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_99_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_99_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1693_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1695_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1697_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1699_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1701_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1703_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1705_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1707_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1709_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1711_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1713_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1715_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1717_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1719_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1721_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1723_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1725_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1727_nl = LOOPK2_and_99_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_47_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_47_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_155_nl, {LOOPK2_LOOPK2_nor_48_nl , LOOPK2_else_and_1693_nl ,
      LOOPK2_else_and_1695_nl , LOOPK2_else_and_1697_nl , LOOPK2_else_and_1699_nl
      , LOOPK2_else_and_1701_nl , LOOPK2_else_and_1703_nl , LOOPK2_else_and_1705_nl
      , LOOPK2_else_and_1707_nl , LOOPK2_else_and_1709_nl , LOOPK2_else_and_1711_nl
      , LOOPK2_else_and_1713_nl , LOOPK2_else_and_1715_nl , LOOPK2_else_and_1717_nl
      , LOOPK2_else_and_1719_nl , LOOPK2_else_and_1721_nl , LOOPK2_else_and_1723_nl
      , LOOPK2_else_and_1725_nl , LOOPK2_else_and_1727_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_538_nl = ~ LOOPK2_and_98_cse_sva_1;
  assign LOOPK2_if_and_154_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_8_lpi_5, LOOPK2_if_not_538_nl);
  assign LOOPK2_LOOPK2_nor_9_nl = ~((~(((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_98_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_98_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_289_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_291_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_293_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_295_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_297_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_299_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_301_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_303_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_305_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_307_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_309_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_311_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_313_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_315_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_317_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_319_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_321_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_323_nl = LOOPK2_and_98_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_8_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_8_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_154_nl, {LOOPK2_LOOPK2_nor_9_nl , LOOPK2_else_and_289_nl , LOOPK2_else_and_291_nl
      , LOOPK2_else_and_293_nl , LOOPK2_else_and_295_nl , LOOPK2_else_and_297_nl
      , LOOPK2_else_and_299_nl , LOOPK2_else_and_301_nl , LOOPK2_else_and_303_nl
      , LOOPK2_else_and_305_nl , LOOPK2_else_and_307_nl , LOOPK2_else_and_309_nl
      , LOOPK2_else_and_311_nl , LOOPK2_else_and_313_nl , LOOPK2_else_and_315_nl
      , LOOPK2_else_and_317_nl , LOOPK2_else_and_319_nl , LOOPK2_else_and_321_nl
      , LOOPK2_else_and_323_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_556_nl = ~ LOOPK2_and_97_cse_sva_1;
  assign LOOPK2_if_and_153_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_46_lpi_5, LOOPK2_if_not_556_nl);
  assign LOOPK2_LOOPK2_nor_47_nl = ~((~(((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_97_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_97_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1657_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1659_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1661_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1663_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1665_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1667_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1669_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1671_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1673_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1675_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1677_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1679_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1681_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1683_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1685_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1687_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1689_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1691_nl = LOOPK2_and_97_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_46_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_46_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_153_nl, {LOOPK2_LOOPK2_nor_47_nl , LOOPK2_else_and_1657_nl ,
      LOOPK2_else_and_1659_nl , LOOPK2_else_and_1661_nl , LOOPK2_else_and_1663_nl
      , LOOPK2_else_and_1665_nl , LOOPK2_else_and_1667_nl , LOOPK2_else_and_1669_nl
      , LOOPK2_else_and_1671_nl , LOOPK2_else_and_1673_nl , LOOPK2_else_and_1675_nl
      , LOOPK2_else_and_1677_nl , LOOPK2_else_and_1679_nl , LOOPK2_else_and_1681_nl
      , LOOPK2_else_and_1683_nl , LOOPK2_else_and_1685_nl , LOOPK2_else_and_1687_nl
      , LOOPK2_else_and_1689_nl , LOOPK2_else_and_1691_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_574_nl = ~ LOOPK2_and_96_cse_sva_1;
  assign LOOPK2_if_and_152_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_9_lpi_5, LOOPK2_if_not_574_nl);
  assign LOOPK2_LOOPK2_nor_10_nl = ~((~(((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_96_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_96_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_325_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_327_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_329_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_331_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_333_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_335_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_337_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_339_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_341_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_343_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_345_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_347_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_349_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_351_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_353_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_355_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_357_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_359_nl = LOOPK2_and_96_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_9_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_9_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_152_nl, {LOOPK2_LOOPK2_nor_10_nl , LOOPK2_else_and_325_nl , LOOPK2_else_and_327_nl
      , LOOPK2_else_and_329_nl , LOOPK2_else_and_331_nl , LOOPK2_else_and_333_nl
      , LOOPK2_else_and_335_nl , LOOPK2_else_and_337_nl , LOOPK2_else_and_339_nl
      , LOOPK2_else_and_341_nl , LOOPK2_else_and_343_nl , LOOPK2_else_and_345_nl
      , LOOPK2_else_and_347_nl , LOOPK2_else_and_349_nl , LOOPK2_else_and_351_nl
      , LOOPK2_else_and_353_nl , LOOPK2_else_and_355_nl , LOOPK2_else_and_357_nl
      , LOOPK2_else_and_359_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_592_nl = ~ LOOPK2_and_95_cse_sva_1;
  assign LOOPK2_if_and_151_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_45_lpi_5, LOOPK2_if_not_592_nl);
  assign LOOPK2_LOOPK2_nor_46_nl = ~((~(((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_95_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_95_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1621_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1623_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1625_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1627_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1629_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1631_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1633_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1635_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1637_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1639_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1641_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1643_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1645_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1647_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1649_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1651_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1653_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1655_nl = LOOPK2_and_95_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_45_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_45_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_151_nl, {LOOPK2_LOOPK2_nor_46_nl , LOOPK2_else_and_1621_nl ,
      LOOPK2_else_and_1623_nl , LOOPK2_else_and_1625_nl , LOOPK2_else_and_1627_nl
      , LOOPK2_else_and_1629_nl , LOOPK2_else_and_1631_nl , LOOPK2_else_and_1633_nl
      , LOOPK2_else_and_1635_nl , LOOPK2_else_and_1637_nl , LOOPK2_else_and_1639_nl
      , LOOPK2_else_and_1641_nl , LOOPK2_else_and_1643_nl , LOOPK2_else_and_1645_nl
      , LOOPK2_else_and_1647_nl , LOOPK2_else_and_1649_nl , LOOPK2_else_and_1651_nl
      , LOOPK2_else_and_1653_nl , LOOPK2_else_and_1655_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_610_nl = ~ LOOPK2_and_94_cse_sva_1;
  assign LOOPK2_if_and_150_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_10_lpi_5, LOOPK2_if_not_610_nl);
  assign LOOPK2_LOOPK2_nor_11_nl = ~((~(((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_94_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_94_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_361_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_363_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_365_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_367_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_369_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_371_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_373_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_375_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_377_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_379_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_381_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_383_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_385_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_387_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_389_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_391_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_393_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_395_nl = LOOPK2_and_94_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_10_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_10_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_150_nl, {LOOPK2_LOOPK2_nor_11_nl , LOOPK2_else_and_361_nl , LOOPK2_else_and_363_nl
      , LOOPK2_else_and_365_nl , LOOPK2_else_and_367_nl , LOOPK2_else_and_369_nl
      , LOOPK2_else_and_371_nl , LOOPK2_else_and_373_nl , LOOPK2_else_and_375_nl
      , LOOPK2_else_and_377_nl , LOOPK2_else_and_379_nl , LOOPK2_else_and_381_nl
      , LOOPK2_else_and_383_nl , LOOPK2_else_and_385_nl , LOOPK2_else_and_387_nl
      , LOOPK2_else_and_389_nl , LOOPK2_else_and_391_nl , LOOPK2_else_and_393_nl
      , LOOPK2_else_and_395_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_628_nl = ~ LOOPK2_and_93_cse_sva_1;
  assign LOOPK2_if_and_149_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_44_lpi_5, LOOPK2_if_not_628_nl);
  assign LOOPK2_LOOPK2_nor_45_nl = ~((~(((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_93_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_93_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1585_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1587_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1589_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1591_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1593_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1595_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1597_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1599_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1601_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1603_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1605_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1607_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1609_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1611_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1613_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1615_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1617_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1619_nl = LOOPK2_and_93_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_44_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_44_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_149_nl, {LOOPK2_LOOPK2_nor_45_nl , LOOPK2_else_and_1585_nl ,
      LOOPK2_else_and_1587_nl , LOOPK2_else_and_1589_nl , LOOPK2_else_and_1591_nl
      , LOOPK2_else_and_1593_nl , LOOPK2_else_and_1595_nl , LOOPK2_else_and_1597_nl
      , LOOPK2_else_and_1599_nl , LOOPK2_else_and_1601_nl , LOOPK2_else_and_1603_nl
      , LOOPK2_else_and_1605_nl , LOOPK2_else_and_1607_nl , LOOPK2_else_and_1609_nl
      , LOOPK2_else_and_1611_nl , LOOPK2_else_and_1613_nl , LOOPK2_else_and_1615_nl
      , LOOPK2_else_and_1617_nl , LOOPK2_else_and_1619_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_646_nl = ~ LOOPK2_and_92_cse_sva_1;
  assign LOOPK2_if_and_148_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_11_lpi_5, LOOPK2_if_not_646_nl);
  assign LOOPK2_LOOPK2_nor_12_nl = ~((~(((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_92_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_92_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_397_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_399_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_401_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_403_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_405_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_407_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_409_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_411_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_413_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_415_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_417_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_419_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_421_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_423_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_425_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_427_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_429_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_431_nl = LOOPK2_and_92_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_11_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_11_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_148_nl, {LOOPK2_LOOPK2_nor_12_nl , LOOPK2_else_and_397_nl , LOOPK2_else_and_399_nl
      , LOOPK2_else_and_401_nl , LOOPK2_else_and_403_nl , LOOPK2_else_and_405_nl
      , LOOPK2_else_and_407_nl , LOOPK2_else_and_409_nl , LOOPK2_else_and_411_nl
      , LOOPK2_else_and_413_nl , LOOPK2_else_and_415_nl , LOOPK2_else_and_417_nl
      , LOOPK2_else_and_419_nl , LOOPK2_else_and_421_nl , LOOPK2_else_and_423_nl
      , LOOPK2_else_and_425_nl , LOOPK2_else_and_427_nl , LOOPK2_else_and_429_nl
      , LOOPK2_else_and_431_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_664_nl = ~ LOOPK2_and_91_cse_sva_1;
  assign LOOPK2_if_and_147_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_43_lpi_5, LOOPK2_if_not_664_nl);
  assign LOOPK2_LOOPK2_nor_44_nl = ~((~(((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_91_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_91_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1549_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1551_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1553_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1555_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1557_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1559_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1561_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1563_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1565_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1567_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1569_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1571_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1573_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1575_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1577_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1579_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1581_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1583_nl = LOOPK2_and_91_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_43_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_43_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_147_nl, {LOOPK2_LOOPK2_nor_44_nl , LOOPK2_else_and_1549_nl ,
      LOOPK2_else_and_1551_nl , LOOPK2_else_and_1553_nl , LOOPK2_else_and_1555_nl
      , LOOPK2_else_and_1557_nl , LOOPK2_else_and_1559_nl , LOOPK2_else_and_1561_nl
      , LOOPK2_else_and_1563_nl , LOOPK2_else_and_1565_nl , LOOPK2_else_and_1567_nl
      , LOOPK2_else_and_1569_nl , LOOPK2_else_and_1571_nl , LOOPK2_else_and_1573_nl
      , LOOPK2_else_and_1575_nl , LOOPK2_else_and_1577_nl , LOOPK2_else_and_1579_nl
      , LOOPK2_else_and_1581_nl , LOOPK2_else_and_1583_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_682_nl = ~ LOOPK2_and_90_cse_sva_1;
  assign LOOPK2_if_and_146_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_12_lpi_5, LOOPK2_if_not_682_nl);
  assign LOOPK2_LOOPK2_nor_13_nl = ~((~(((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_90_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_90_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_433_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_435_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_437_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_439_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_441_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_443_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_445_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_447_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_449_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_451_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_453_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_455_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_457_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_459_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_461_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_463_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_465_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_467_nl = LOOPK2_and_90_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_12_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_12_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_146_nl, {LOOPK2_LOOPK2_nor_13_nl , LOOPK2_else_and_433_nl , LOOPK2_else_and_435_nl
      , LOOPK2_else_and_437_nl , LOOPK2_else_and_439_nl , LOOPK2_else_and_441_nl
      , LOOPK2_else_and_443_nl , LOOPK2_else_and_445_nl , LOOPK2_else_and_447_nl
      , LOOPK2_else_and_449_nl , LOOPK2_else_and_451_nl , LOOPK2_else_and_453_nl
      , LOOPK2_else_and_455_nl , LOOPK2_else_and_457_nl , LOOPK2_else_and_459_nl
      , LOOPK2_else_and_461_nl , LOOPK2_else_and_463_nl , LOOPK2_else_and_465_nl
      , LOOPK2_else_and_467_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_700_nl = ~ LOOPK2_and_89_cse_sva_1;
  assign LOOPK2_if_and_145_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_42_lpi_5, LOOPK2_if_not_700_nl);
  assign LOOPK2_LOOPK2_nor_43_nl = ~((~(((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_89_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_89_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1513_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1515_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1517_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1519_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1521_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1523_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1525_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1527_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1529_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1531_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1533_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1535_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1537_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1539_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1541_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1543_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1545_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1547_nl = LOOPK2_and_89_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_42_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_42_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_145_nl, {LOOPK2_LOOPK2_nor_43_nl , LOOPK2_else_and_1513_nl ,
      LOOPK2_else_and_1515_nl , LOOPK2_else_and_1517_nl , LOOPK2_else_and_1519_nl
      , LOOPK2_else_and_1521_nl , LOOPK2_else_and_1523_nl , LOOPK2_else_and_1525_nl
      , LOOPK2_else_and_1527_nl , LOOPK2_else_and_1529_nl , LOOPK2_else_and_1531_nl
      , LOOPK2_else_and_1533_nl , LOOPK2_else_and_1535_nl , LOOPK2_else_and_1537_nl
      , LOOPK2_else_and_1539_nl , LOOPK2_else_and_1541_nl , LOOPK2_else_and_1543_nl
      , LOOPK2_else_and_1545_nl , LOOPK2_else_and_1547_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_718_nl = ~ LOOPK2_and_88_cse_sva_1;
  assign LOOPK2_if_and_144_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_13_lpi_5, LOOPK2_if_not_718_nl);
  assign LOOPK2_LOOPK2_nor_14_nl = ~((~(((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_88_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_88_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_469_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_471_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_473_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_475_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_477_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_479_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_481_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_483_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_485_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_487_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_489_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_491_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_493_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_495_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_497_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_499_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_501_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_503_nl = LOOPK2_and_88_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_13_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_13_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_144_nl, {LOOPK2_LOOPK2_nor_14_nl , LOOPK2_else_and_469_nl , LOOPK2_else_and_471_nl
      , LOOPK2_else_and_473_nl , LOOPK2_else_and_475_nl , LOOPK2_else_and_477_nl
      , LOOPK2_else_and_479_nl , LOOPK2_else_and_481_nl , LOOPK2_else_and_483_nl
      , LOOPK2_else_and_485_nl , LOOPK2_else_and_487_nl , LOOPK2_else_and_489_nl
      , LOOPK2_else_and_491_nl , LOOPK2_else_and_493_nl , LOOPK2_else_and_495_nl
      , LOOPK2_else_and_497_nl , LOOPK2_else_and_499_nl , LOOPK2_else_and_501_nl
      , LOOPK2_else_and_503_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_736_nl = ~ LOOPK2_and_87_cse_sva_1;
  assign LOOPK2_if_and_143_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_41_lpi_5, LOOPK2_if_not_736_nl);
  assign LOOPK2_LOOPK2_nor_42_nl = ~((~(((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_87_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_87_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1477_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1479_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1481_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1483_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1485_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1487_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1489_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1491_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1493_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1495_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1497_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1499_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1501_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1503_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1505_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1507_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1509_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1511_nl = LOOPK2_and_87_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_41_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_41_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_143_nl, {LOOPK2_LOOPK2_nor_42_nl , LOOPK2_else_and_1477_nl ,
      LOOPK2_else_and_1479_nl , LOOPK2_else_and_1481_nl , LOOPK2_else_and_1483_nl
      , LOOPK2_else_and_1485_nl , LOOPK2_else_and_1487_nl , LOOPK2_else_and_1489_nl
      , LOOPK2_else_and_1491_nl , LOOPK2_else_and_1493_nl , LOOPK2_else_and_1495_nl
      , LOOPK2_else_and_1497_nl , LOOPK2_else_and_1499_nl , LOOPK2_else_and_1501_nl
      , LOOPK2_else_and_1503_nl , LOOPK2_else_and_1505_nl , LOOPK2_else_and_1507_nl
      , LOOPK2_else_and_1509_nl , LOOPK2_else_and_1511_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_754_nl = ~ LOOPK2_and_86_cse_sva_1;
  assign LOOPK2_if_and_142_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_14_lpi_5, LOOPK2_if_not_754_nl);
  assign LOOPK2_LOOPK2_nor_15_nl = ~((~(((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_86_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_86_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_505_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_507_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_509_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_511_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_513_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_515_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_517_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_519_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_521_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_523_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_525_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_527_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_529_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_531_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_533_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_535_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_537_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_539_nl = LOOPK2_and_86_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_14_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_14_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_142_nl, {LOOPK2_LOOPK2_nor_15_nl , LOOPK2_else_and_505_nl , LOOPK2_else_and_507_nl
      , LOOPK2_else_and_509_nl , LOOPK2_else_and_511_nl , LOOPK2_else_and_513_nl
      , LOOPK2_else_and_515_nl , LOOPK2_else_and_517_nl , LOOPK2_else_and_519_nl
      , LOOPK2_else_and_521_nl , LOOPK2_else_and_523_nl , LOOPK2_else_and_525_nl
      , LOOPK2_else_and_527_nl , LOOPK2_else_and_529_nl , LOOPK2_else_and_531_nl
      , LOOPK2_else_and_533_nl , LOOPK2_else_and_535_nl , LOOPK2_else_and_537_nl
      , LOOPK2_else_and_539_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_772_nl = ~ LOOPK2_and_85_cse_sva_1;
  assign LOOPK2_if_and_141_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_40_lpi_5, LOOPK2_if_not_772_nl);
  assign LOOPK2_LOOPK2_nor_41_nl = ~((~(((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_85_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_85_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1441_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1443_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1445_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1447_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1449_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1451_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1453_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1455_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1457_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1459_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1461_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1463_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1465_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1467_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1469_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1471_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1473_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1475_nl = LOOPK2_and_85_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_40_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_40_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_141_nl, {LOOPK2_LOOPK2_nor_41_nl , LOOPK2_else_and_1441_nl ,
      LOOPK2_else_and_1443_nl , LOOPK2_else_and_1445_nl , LOOPK2_else_and_1447_nl
      , LOOPK2_else_and_1449_nl , LOOPK2_else_and_1451_nl , LOOPK2_else_and_1453_nl
      , LOOPK2_else_and_1455_nl , LOOPK2_else_and_1457_nl , LOOPK2_else_and_1459_nl
      , LOOPK2_else_and_1461_nl , LOOPK2_else_and_1463_nl , LOOPK2_else_and_1465_nl
      , LOOPK2_else_and_1467_nl , LOOPK2_else_and_1469_nl , LOOPK2_else_and_1471_nl
      , LOOPK2_else_and_1473_nl , LOOPK2_else_and_1475_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_790_nl = ~ LOOPK2_and_84_cse_sva_1;
  assign LOOPK2_if_and_140_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_15_lpi_5, LOOPK2_if_not_790_nl);
  assign LOOPK2_LOOPK2_nor_16_nl = ~((~(((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_84_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_84_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_541_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_543_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_545_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_547_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_549_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_551_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_553_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_555_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_557_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_559_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_561_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_563_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_565_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_567_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_569_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_571_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_573_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_575_nl = LOOPK2_and_84_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_15_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_15_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_140_nl, {LOOPK2_LOOPK2_nor_16_nl , LOOPK2_else_and_541_nl , LOOPK2_else_and_543_nl
      , LOOPK2_else_and_545_nl , LOOPK2_else_and_547_nl , LOOPK2_else_and_549_nl
      , LOOPK2_else_and_551_nl , LOOPK2_else_and_553_nl , LOOPK2_else_and_555_nl
      , LOOPK2_else_and_557_nl , LOOPK2_else_and_559_nl , LOOPK2_else_and_561_nl
      , LOOPK2_else_and_563_nl , LOOPK2_else_and_565_nl , LOOPK2_else_and_567_nl
      , LOOPK2_else_and_569_nl , LOOPK2_else_and_571_nl , LOOPK2_else_and_573_nl
      , LOOPK2_else_and_575_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_808_nl = ~ LOOPK2_and_83_cse_sva_1;
  assign LOOPK2_if_and_139_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_39_lpi_5, LOOPK2_if_not_808_nl);
  assign LOOPK2_LOOPK2_nor_40_nl = ~((~(((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_83_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_83_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1405_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1407_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1409_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1411_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1413_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1415_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1417_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1419_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1421_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1423_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1425_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1427_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1429_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1431_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1433_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1435_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1437_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1439_nl = LOOPK2_and_83_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_39_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_39_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_139_nl, {LOOPK2_LOOPK2_nor_40_nl , LOOPK2_else_and_1405_nl ,
      LOOPK2_else_and_1407_nl , LOOPK2_else_and_1409_nl , LOOPK2_else_and_1411_nl
      , LOOPK2_else_and_1413_nl , LOOPK2_else_and_1415_nl , LOOPK2_else_and_1417_nl
      , LOOPK2_else_and_1419_nl , LOOPK2_else_and_1421_nl , LOOPK2_else_and_1423_nl
      , LOOPK2_else_and_1425_nl , LOOPK2_else_and_1427_nl , LOOPK2_else_and_1429_nl
      , LOOPK2_else_and_1431_nl , LOOPK2_else_and_1433_nl , LOOPK2_else_and_1435_nl
      , LOOPK2_else_and_1437_nl , LOOPK2_else_and_1439_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_826_nl = ~ LOOPK2_and_82_cse_sva_1;
  assign LOOPK2_if_and_138_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_16_lpi_5, LOOPK2_if_not_826_nl);
  assign LOOPK2_LOOPK2_nor_17_nl = ~((~(((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_82_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_82_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_577_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_579_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_581_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_583_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_585_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_587_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_589_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_591_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_593_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_595_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_597_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_599_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_601_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_603_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_605_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_607_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_609_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_611_nl = LOOPK2_and_82_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_16_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_16_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_138_nl, {LOOPK2_LOOPK2_nor_17_nl , LOOPK2_else_and_577_nl , LOOPK2_else_and_579_nl
      , LOOPK2_else_and_581_nl , LOOPK2_else_and_583_nl , LOOPK2_else_and_585_nl
      , LOOPK2_else_and_587_nl , LOOPK2_else_and_589_nl , LOOPK2_else_and_591_nl
      , LOOPK2_else_and_593_nl , LOOPK2_else_and_595_nl , LOOPK2_else_and_597_nl
      , LOOPK2_else_and_599_nl , LOOPK2_else_and_601_nl , LOOPK2_else_and_603_nl
      , LOOPK2_else_and_605_nl , LOOPK2_else_and_607_nl , LOOPK2_else_and_609_nl
      , LOOPK2_else_and_611_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_844_nl = ~ LOOPK2_and_81_cse_sva_1;
  assign LOOPK2_if_and_137_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_38_lpi_5, LOOPK2_if_not_844_nl);
  assign LOOPK2_LOOPK2_nor_39_nl = ~((~(((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_81_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_81_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1369_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1371_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1373_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1375_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1377_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1379_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1381_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1383_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1385_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1387_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1389_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1391_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1393_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1395_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1397_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1399_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1401_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1403_nl = LOOPK2_and_81_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_38_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_38_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_137_nl, {LOOPK2_LOOPK2_nor_39_nl , LOOPK2_else_and_1369_nl ,
      LOOPK2_else_and_1371_nl , LOOPK2_else_and_1373_nl , LOOPK2_else_and_1375_nl
      , LOOPK2_else_and_1377_nl , LOOPK2_else_and_1379_nl , LOOPK2_else_and_1381_nl
      , LOOPK2_else_and_1383_nl , LOOPK2_else_and_1385_nl , LOOPK2_else_and_1387_nl
      , LOOPK2_else_and_1389_nl , LOOPK2_else_and_1391_nl , LOOPK2_else_and_1393_nl
      , LOOPK2_else_and_1395_nl , LOOPK2_else_and_1397_nl , LOOPK2_else_and_1399_nl
      , LOOPK2_else_and_1401_nl , LOOPK2_else_and_1403_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_862_nl = ~ LOOPK2_and_80_cse_sva_1;
  assign LOOPK2_if_and_136_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_17_lpi_5, LOOPK2_if_not_862_nl);
  assign LOOPK2_LOOPK2_nor_18_nl = ~((~(((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_80_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_80_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_613_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_615_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_617_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_619_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_621_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_623_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_625_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_627_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_629_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_631_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_633_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_635_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_637_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_639_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_641_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_643_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_645_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_647_nl = LOOPK2_and_80_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_17_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_17_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_136_nl, {LOOPK2_LOOPK2_nor_18_nl , LOOPK2_else_and_613_nl , LOOPK2_else_and_615_nl
      , LOOPK2_else_and_617_nl , LOOPK2_else_and_619_nl , LOOPK2_else_and_621_nl
      , LOOPK2_else_and_623_nl , LOOPK2_else_and_625_nl , LOOPK2_else_and_627_nl
      , LOOPK2_else_and_629_nl , LOOPK2_else_and_631_nl , LOOPK2_else_and_633_nl
      , LOOPK2_else_and_635_nl , LOOPK2_else_and_637_nl , LOOPK2_else_and_639_nl
      , LOOPK2_else_and_641_nl , LOOPK2_else_and_643_nl , LOOPK2_else_and_645_nl
      , LOOPK2_else_and_647_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_880_nl = ~ LOOPK2_and_79_cse_sva_1;
  assign LOOPK2_if_and_135_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_37_lpi_5, LOOPK2_if_not_880_nl);
  assign LOOPK2_LOOPK2_nor_38_nl = ~((~(((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_79_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_79_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1333_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1335_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1337_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1339_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1341_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1343_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1345_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1347_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1349_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1351_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1353_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1355_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1357_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1359_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1361_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1363_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1365_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1367_nl = LOOPK2_and_79_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_37_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_37_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_135_nl, {LOOPK2_LOOPK2_nor_38_nl , LOOPK2_else_and_1333_nl ,
      LOOPK2_else_and_1335_nl , LOOPK2_else_and_1337_nl , LOOPK2_else_and_1339_nl
      , LOOPK2_else_and_1341_nl , LOOPK2_else_and_1343_nl , LOOPK2_else_and_1345_nl
      , LOOPK2_else_and_1347_nl , LOOPK2_else_and_1349_nl , LOOPK2_else_and_1351_nl
      , LOOPK2_else_and_1353_nl , LOOPK2_else_and_1355_nl , LOOPK2_else_and_1357_nl
      , LOOPK2_else_and_1359_nl , LOOPK2_else_and_1361_nl , LOOPK2_else_and_1363_nl
      , LOOPK2_else_and_1365_nl , LOOPK2_else_and_1367_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_898_nl = ~ LOOPK2_and_78_cse_sva_1;
  assign LOOPK2_if_and_134_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_18_lpi_5, LOOPK2_if_not_898_nl);
  assign LOOPK2_LOOPK2_nor_19_nl = ~((~(((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_78_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_78_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_649_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_651_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_653_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_655_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_657_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_659_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_661_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_663_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_665_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_667_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_669_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_671_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_673_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_675_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_677_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_679_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_681_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_683_nl = LOOPK2_and_78_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_18_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_18_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_134_nl, {LOOPK2_LOOPK2_nor_19_nl , LOOPK2_else_and_649_nl , LOOPK2_else_and_651_nl
      , LOOPK2_else_and_653_nl , LOOPK2_else_and_655_nl , LOOPK2_else_and_657_nl
      , LOOPK2_else_and_659_nl , LOOPK2_else_and_661_nl , LOOPK2_else_and_663_nl
      , LOOPK2_else_and_665_nl , LOOPK2_else_and_667_nl , LOOPK2_else_and_669_nl
      , LOOPK2_else_and_671_nl , LOOPK2_else_and_673_nl , LOOPK2_else_and_675_nl
      , LOOPK2_else_and_677_nl , LOOPK2_else_and_679_nl , LOOPK2_else_and_681_nl
      , LOOPK2_else_and_683_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_916_nl = ~ LOOPK2_and_77_cse_sva_1;
  assign LOOPK2_if_and_133_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_36_lpi_5, LOOPK2_if_not_916_nl);
  assign LOOPK2_LOOPK2_nor_37_nl = ~((~(((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_77_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_77_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1297_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1299_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1301_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1303_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1305_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1307_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1309_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1311_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1313_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1315_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1317_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1319_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1321_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1323_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1325_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1327_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1329_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1331_nl = LOOPK2_and_77_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_36_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_36_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_133_nl, {LOOPK2_LOOPK2_nor_37_nl , LOOPK2_else_and_1297_nl ,
      LOOPK2_else_and_1299_nl , LOOPK2_else_and_1301_nl , LOOPK2_else_and_1303_nl
      , LOOPK2_else_and_1305_nl , LOOPK2_else_and_1307_nl , LOOPK2_else_and_1309_nl
      , LOOPK2_else_and_1311_nl , LOOPK2_else_and_1313_nl , LOOPK2_else_and_1315_nl
      , LOOPK2_else_and_1317_nl , LOOPK2_else_and_1319_nl , LOOPK2_else_and_1321_nl
      , LOOPK2_else_and_1323_nl , LOOPK2_else_and_1325_nl , LOOPK2_else_and_1327_nl
      , LOOPK2_else_and_1329_nl , LOOPK2_else_and_1331_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_934_nl = ~ LOOPK2_and_76_cse_sva_1;
  assign LOOPK2_if_and_132_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_19_lpi_5, LOOPK2_if_not_934_nl);
  assign LOOPK2_LOOPK2_nor_20_nl = ~((~(((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_76_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_76_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_685_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_687_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_689_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_691_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_693_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_695_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_697_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_699_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_701_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_703_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_705_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_707_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_709_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_711_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_713_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_715_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_717_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_719_nl = LOOPK2_and_76_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_19_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_19_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_132_nl, {LOOPK2_LOOPK2_nor_20_nl , LOOPK2_else_and_685_nl , LOOPK2_else_and_687_nl
      , LOOPK2_else_and_689_nl , LOOPK2_else_and_691_nl , LOOPK2_else_and_693_nl
      , LOOPK2_else_and_695_nl , LOOPK2_else_and_697_nl , LOOPK2_else_and_699_nl
      , LOOPK2_else_and_701_nl , LOOPK2_else_and_703_nl , LOOPK2_else_and_705_nl
      , LOOPK2_else_and_707_nl , LOOPK2_else_and_709_nl , LOOPK2_else_and_711_nl
      , LOOPK2_else_and_713_nl , LOOPK2_else_and_715_nl , LOOPK2_else_and_717_nl
      , LOOPK2_else_and_719_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_952_nl = ~ LOOPK2_and_75_cse_sva_1;
  assign LOOPK2_if_and_131_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_35_lpi_5, LOOPK2_if_not_952_nl);
  assign LOOPK2_LOOPK2_nor_36_nl = ~((~(((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_75_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_75_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1261_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1263_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1265_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1267_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1269_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1271_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1273_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1275_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1277_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1279_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1281_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1283_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1285_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1287_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1289_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1291_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1293_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1295_nl = LOOPK2_and_75_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_35_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_35_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_131_nl, {LOOPK2_LOOPK2_nor_36_nl , LOOPK2_else_and_1261_nl ,
      LOOPK2_else_and_1263_nl , LOOPK2_else_and_1265_nl , LOOPK2_else_and_1267_nl
      , LOOPK2_else_and_1269_nl , LOOPK2_else_and_1271_nl , LOOPK2_else_and_1273_nl
      , LOOPK2_else_and_1275_nl , LOOPK2_else_and_1277_nl , LOOPK2_else_and_1279_nl
      , LOOPK2_else_and_1281_nl , LOOPK2_else_and_1283_nl , LOOPK2_else_and_1285_nl
      , LOOPK2_else_and_1287_nl , LOOPK2_else_and_1289_nl , LOOPK2_else_and_1291_nl
      , LOOPK2_else_and_1293_nl , LOOPK2_else_and_1295_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_970_nl = ~ LOOPK2_and_74_cse_sva_1;
  assign LOOPK2_if_and_130_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_20_lpi_5, LOOPK2_if_not_970_nl);
  assign LOOPK2_LOOPK2_nor_21_nl = ~((~(((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_74_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_74_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_721_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_723_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_725_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_727_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_729_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_731_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_733_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_735_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_737_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_739_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_741_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_743_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_745_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_747_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_749_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_751_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_753_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_755_nl = LOOPK2_and_74_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_20_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_20_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_130_nl, {LOOPK2_LOOPK2_nor_21_nl , LOOPK2_else_and_721_nl , LOOPK2_else_and_723_nl
      , LOOPK2_else_and_725_nl , LOOPK2_else_and_727_nl , LOOPK2_else_and_729_nl
      , LOOPK2_else_and_731_nl , LOOPK2_else_and_733_nl , LOOPK2_else_and_735_nl
      , LOOPK2_else_and_737_nl , LOOPK2_else_and_739_nl , LOOPK2_else_and_741_nl
      , LOOPK2_else_and_743_nl , LOOPK2_else_and_745_nl , LOOPK2_else_and_747_nl
      , LOOPK2_else_and_749_nl , LOOPK2_else_and_751_nl , LOOPK2_else_and_753_nl
      , LOOPK2_else_and_755_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_988_nl = ~ LOOPK2_and_73_cse_sva_1;
  assign LOOPK2_if_and_129_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_34_lpi_5, LOOPK2_if_not_988_nl);
  assign LOOPK2_LOOPK2_nor_35_nl = ~((~(((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_73_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_73_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1225_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1227_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1229_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1231_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1233_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1235_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1237_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1239_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1241_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1243_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1245_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1247_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1249_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1251_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1253_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1255_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1257_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1259_nl = LOOPK2_and_73_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_34_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_34_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_129_nl, {LOOPK2_LOOPK2_nor_35_nl , LOOPK2_else_and_1225_nl ,
      LOOPK2_else_and_1227_nl , LOOPK2_else_and_1229_nl , LOOPK2_else_and_1231_nl
      , LOOPK2_else_and_1233_nl , LOOPK2_else_and_1235_nl , LOOPK2_else_and_1237_nl
      , LOOPK2_else_and_1239_nl , LOOPK2_else_and_1241_nl , LOOPK2_else_and_1243_nl
      , LOOPK2_else_and_1245_nl , LOOPK2_else_and_1247_nl , LOOPK2_else_and_1249_nl
      , LOOPK2_else_and_1251_nl , LOOPK2_else_and_1253_nl , LOOPK2_else_and_1255_nl
      , LOOPK2_else_and_1257_nl , LOOPK2_else_and_1259_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1006_nl = ~ LOOPK2_and_72_cse_sva_1;
  assign LOOPK2_if_and_128_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_21_lpi_5, LOOPK2_if_not_1006_nl);
  assign LOOPK2_LOOPK2_nor_22_nl = ~((~(((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_72_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_72_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_757_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_759_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_761_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_763_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_765_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_767_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_769_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_771_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_773_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_775_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_777_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_779_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_781_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_783_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_785_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_787_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_789_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_791_nl = LOOPK2_and_72_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_21_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_21_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_128_nl, {LOOPK2_LOOPK2_nor_22_nl , LOOPK2_else_and_757_nl , LOOPK2_else_and_759_nl
      , LOOPK2_else_and_761_nl , LOOPK2_else_and_763_nl , LOOPK2_else_and_765_nl
      , LOOPK2_else_and_767_nl , LOOPK2_else_and_769_nl , LOOPK2_else_and_771_nl
      , LOOPK2_else_and_773_nl , LOOPK2_else_and_775_nl , LOOPK2_else_and_777_nl
      , LOOPK2_else_and_779_nl , LOOPK2_else_and_781_nl , LOOPK2_else_and_783_nl
      , LOOPK2_else_and_785_nl , LOOPK2_else_and_787_nl , LOOPK2_else_and_789_nl
      , LOOPK2_else_and_791_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1024_nl = ~ LOOPK2_and_71_cse_sva_1;
  assign LOOPK2_if_and_127_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_33_lpi_5, LOOPK2_if_not_1024_nl);
  assign LOOPK2_LOOPK2_nor_34_nl = ~((~(((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_71_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_71_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1189_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1191_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1193_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1195_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1197_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1199_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1201_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1203_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1205_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1207_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1209_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1211_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1213_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1215_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1217_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1219_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1221_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1223_nl = LOOPK2_and_71_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_33_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_33_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_127_nl, {LOOPK2_LOOPK2_nor_34_nl , LOOPK2_else_and_1189_nl ,
      LOOPK2_else_and_1191_nl , LOOPK2_else_and_1193_nl , LOOPK2_else_and_1195_nl
      , LOOPK2_else_and_1197_nl , LOOPK2_else_and_1199_nl , LOOPK2_else_and_1201_nl
      , LOOPK2_else_and_1203_nl , LOOPK2_else_and_1205_nl , LOOPK2_else_and_1207_nl
      , LOOPK2_else_and_1209_nl , LOOPK2_else_and_1211_nl , LOOPK2_else_and_1213_nl
      , LOOPK2_else_and_1215_nl , LOOPK2_else_and_1217_nl , LOOPK2_else_and_1219_nl
      , LOOPK2_else_and_1221_nl , LOOPK2_else_and_1223_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1042_nl = ~ LOOPK2_and_70_cse_sva_1;
  assign LOOPK2_if_and_126_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_22_lpi_5, LOOPK2_if_not_1042_nl);
  assign LOOPK2_LOOPK2_nor_23_nl = ~((~(((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_70_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_70_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_793_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_795_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_797_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_799_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_801_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_803_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_805_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_807_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_809_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_811_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_813_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_815_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_817_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_819_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_821_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_823_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_825_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_827_nl = LOOPK2_and_70_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_22_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_22_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_126_nl, {LOOPK2_LOOPK2_nor_23_nl , LOOPK2_else_and_793_nl , LOOPK2_else_and_795_nl
      , LOOPK2_else_and_797_nl , LOOPK2_else_and_799_nl , LOOPK2_else_and_801_nl
      , LOOPK2_else_and_803_nl , LOOPK2_else_and_805_nl , LOOPK2_else_and_807_nl
      , LOOPK2_else_and_809_nl , LOOPK2_else_and_811_nl , LOOPK2_else_and_813_nl
      , LOOPK2_else_and_815_nl , LOOPK2_else_and_817_nl , LOOPK2_else_and_819_nl
      , LOOPK2_else_and_821_nl , LOOPK2_else_and_823_nl , LOOPK2_else_and_825_nl
      , LOOPK2_else_and_827_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1060_nl = ~ LOOPK2_and_69_cse_sva_1;
  assign LOOPK2_if_and_125_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_32_lpi_5, LOOPK2_if_not_1060_nl);
  assign LOOPK2_LOOPK2_nor_33_nl = ~((~(((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_69_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_69_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1153_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1155_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1157_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1159_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1161_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1163_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1165_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1167_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1169_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1171_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1173_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1175_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1177_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1179_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1181_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1183_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1185_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1187_nl = LOOPK2_and_69_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_32_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_32_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_125_nl, {LOOPK2_LOOPK2_nor_33_nl , LOOPK2_else_and_1153_nl ,
      LOOPK2_else_and_1155_nl , LOOPK2_else_and_1157_nl , LOOPK2_else_and_1159_nl
      , LOOPK2_else_and_1161_nl , LOOPK2_else_and_1163_nl , LOOPK2_else_and_1165_nl
      , LOOPK2_else_and_1167_nl , LOOPK2_else_and_1169_nl , LOOPK2_else_and_1171_nl
      , LOOPK2_else_and_1173_nl , LOOPK2_else_and_1175_nl , LOOPK2_else_and_1177_nl
      , LOOPK2_else_and_1179_nl , LOOPK2_else_and_1181_nl , LOOPK2_else_and_1183_nl
      , LOOPK2_else_and_1185_nl , LOOPK2_else_and_1187_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1078_nl = ~ LOOPK2_and_68_cse_sva_1;
  assign LOOPK2_if_and_124_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_23_lpi_5, LOOPK2_if_not_1078_nl);
  assign LOOPK2_LOOPK2_nor_24_nl = ~((~(((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_68_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_68_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_829_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_831_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_833_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_835_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_837_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_839_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_841_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_843_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_845_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_847_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_849_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_851_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_853_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_855_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_857_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_859_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_861_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_863_nl = LOOPK2_and_68_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_23_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_23_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_124_nl, {LOOPK2_LOOPK2_nor_24_nl , LOOPK2_else_and_829_nl , LOOPK2_else_and_831_nl
      , LOOPK2_else_and_833_nl , LOOPK2_else_and_835_nl , LOOPK2_else_and_837_nl
      , LOOPK2_else_and_839_nl , LOOPK2_else_and_841_nl , LOOPK2_else_and_843_nl
      , LOOPK2_else_and_845_nl , LOOPK2_else_and_847_nl , LOOPK2_else_and_849_nl
      , LOOPK2_else_and_851_nl , LOOPK2_else_and_853_nl , LOOPK2_else_and_855_nl
      , LOOPK2_else_and_857_nl , LOOPK2_else_and_859_nl , LOOPK2_else_and_861_nl
      , LOOPK2_else_and_863_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1096_nl = ~ LOOPK2_and_67_cse_sva_1;
  assign LOOPK2_if_and_123_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_31_lpi_5, LOOPK2_if_not_1096_nl);
  assign LOOPK2_LOOPK2_nor_32_nl = ~((~(((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_67_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_67_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1117_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1119_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1121_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1123_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1125_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1127_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1129_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1131_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1133_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1135_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1137_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1139_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1141_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1143_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1145_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1147_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1149_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1151_nl = LOOPK2_and_67_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_31_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_31_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_123_nl, {LOOPK2_LOOPK2_nor_32_nl , LOOPK2_else_and_1117_nl ,
      LOOPK2_else_and_1119_nl , LOOPK2_else_and_1121_nl , LOOPK2_else_and_1123_nl
      , LOOPK2_else_and_1125_nl , LOOPK2_else_and_1127_nl , LOOPK2_else_and_1129_nl
      , LOOPK2_else_and_1131_nl , LOOPK2_else_and_1133_nl , LOOPK2_else_and_1135_nl
      , LOOPK2_else_and_1137_nl , LOOPK2_else_and_1139_nl , LOOPK2_else_and_1141_nl
      , LOOPK2_else_and_1143_nl , LOOPK2_else_and_1145_nl , LOOPK2_else_and_1147_nl
      , LOOPK2_else_and_1149_nl , LOOPK2_else_and_1151_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1114_nl = ~ LOOPK2_and_66_cse_sva_1;
  assign LOOPK2_if_and_122_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_24_lpi_5, LOOPK2_if_not_1114_nl);
  assign LOOPK2_LOOPK2_nor_25_nl = ~((~(((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_66_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_66_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_865_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_867_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_869_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_871_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_873_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_875_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_877_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_879_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_881_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_883_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_885_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_887_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_889_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_891_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_893_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_895_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_897_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_899_nl = LOOPK2_and_66_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_24_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_24_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_122_nl, {LOOPK2_LOOPK2_nor_25_nl , LOOPK2_else_and_865_nl , LOOPK2_else_and_867_nl
      , LOOPK2_else_and_869_nl , LOOPK2_else_and_871_nl , LOOPK2_else_and_873_nl
      , LOOPK2_else_and_875_nl , LOOPK2_else_and_877_nl , LOOPK2_else_and_879_nl
      , LOOPK2_else_and_881_nl , LOOPK2_else_and_883_nl , LOOPK2_else_and_885_nl
      , LOOPK2_else_and_887_nl , LOOPK2_else_and_889_nl , LOOPK2_else_and_891_nl
      , LOOPK2_else_and_893_nl , LOOPK2_else_and_895_nl , LOOPK2_else_and_897_nl
      , LOOPK2_else_and_899_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1132_nl = ~ LOOPK2_and_65_cse_sva_1;
  assign LOOPK2_if_and_121_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_30_lpi_5, LOOPK2_if_not_1132_nl);
  assign LOOPK2_LOOPK2_nor_31_nl = ~((~(((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_65_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_65_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1081_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1083_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1085_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1087_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1089_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1091_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1093_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1095_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1097_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1099_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1101_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1103_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1105_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1107_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1109_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1111_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1113_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1115_nl = LOOPK2_and_65_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_30_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_30_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_121_nl, {LOOPK2_LOOPK2_nor_31_nl , LOOPK2_else_and_1081_nl ,
      LOOPK2_else_and_1083_nl , LOOPK2_else_and_1085_nl , LOOPK2_else_and_1087_nl
      , LOOPK2_else_and_1089_nl , LOOPK2_else_and_1091_nl , LOOPK2_else_and_1093_nl
      , LOOPK2_else_and_1095_nl , LOOPK2_else_and_1097_nl , LOOPK2_else_and_1099_nl
      , LOOPK2_else_and_1101_nl , LOOPK2_else_and_1103_nl , LOOPK2_else_and_1105_nl
      , LOOPK2_else_and_1107_nl , LOOPK2_else_and_1109_nl , LOOPK2_else_and_1111_nl
      , LOOPK2_else_and_1113_nl , LOOPK2_else_and_1115_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1150_nl = ~ LOOPK2_and_64_cse_sva_1;
  assign LOOPK2_if_and_120_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_25_lpi_5, LOOPK2_if_not_1150_nl);
  assign LOOPK2_LOOPK2_nor_26_nl = ~((~(((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_64_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_64_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_901_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_903_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_905_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_907_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_909_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_911_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_913_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_915_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_917_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_919_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_921_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_923_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_925_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_927_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_929_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_931_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_933_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_935_nl = LOOPK2_and_64_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_25_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_25_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_120_nl, {LOOPK2_LOOPK2_nor_26_nl , LOOPK2_else_and_901_nl , LOOPK2_else_and_903_nl
      , LOOPK2_else_and_905_nl , LOOPK2_else_and_907_nl , LOOPK2_else_and_909_nl
      , LOOPK2_else_and_911_nl , LOOPK2_else_and_913_nl , LOOPK2_else_and_915_nl
      , LOOPK2_else_and_917_nl , LOOPK2_else_and_919_nl , LOOPK2_else_and_921_nl
      , LOOPK2_else_and_923_nl , LOOPK2_else_and_925_nl , LOOPK2_else_and_927_nl
      , LOOPK2_else_and_929_nl , LOOPK2_else_and_931_nl , LOOPK2_else_and_933_nl
      , LOOPK2_else_and_935_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1168_nl = ~ LOOPK2_and_63_cse_sva_1;
  assign LOOPK2_if_and_119_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_29_lpi_5, LOOPK2_if_not_1168_nl);
  assign LOOPK2_LOOPK2_nor_30_nl = ~((~(((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_63_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_63_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1045_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1047_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1049_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1051_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1053_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1055_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1057_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1059_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1061_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1063_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1065_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1067_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1069_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1071_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1073_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1075_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1077_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1079_nl = LOOPK2_and_63_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_29_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_29_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_119_nl, {LOOPK2_LOOPK2_nor_30_nl , LOOPK2_else_and_1045_nl ,
      LOOPK2_else_and_1047_nl , LOOPK2_else_and_1049_nl , LOOPK2_else_and_1051_nl
      , LOOPK2_else_and_1053_nl , LOOPK2_else_and_1055_nl , LOOPK2_else_and_1057_nl
      , LOOPK2_else_and_1059_nl , LOOPK2_else_and_1061_nl , LOOPK2_else_and_1063_nl
      , LOOPK2_else_and_1065_nl , LOOPK2_else_and_1067_nl , LOOPK2_else_and_1069_nl
      , LOOPK2_else_and_1071_nl , LOOPK2_else_and_1073_nl , LOOPK2_else_and_1075_nl
      , LOOPK2_else_and_1077_nl , LOOPK2_else_and_1079_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1186_nl = ~ LOOPK2_and_62_cse_sva_1;
  assign LOOPK2_if_and_118_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_26_lpi_5, LOOPK2_if_not_1186_nl);
  assign LOOPK2_LOOPK2_nor_27_nl = ~((~(((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_62_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_62_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_937_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_939_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_941_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_943_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_945_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_947_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_949_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_951_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_953_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_955_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_957_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_959_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_961_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_963_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_965_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_967_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_969_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_971_nl = LOOPK2_and_62_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_26_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_26_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_118_nl, {LOOPK2_LOOPK2_nor_27_nl , LOOPK2_else_and_937_nl , LOOPK2_else_and_939_nl
      , LOOPK2_else_and_941_nl , LOOPK2_else_and_943_nl , LOOPK2_else_and_945_nl
      , LOOPK2_else_and_947_nl , LOOPK2_else_and_949_nl , LOOPK2_else_and_951_nl
      , LOOPK2_else_and_953_nl , LOOPK2_else_and_955_nl , LOOPK2_else_and_957_nl
      , LOOPK2_else_and_959_nl , LOOPK2_else_and_961_nl , LOOPK2_else_and_963_nl
      , LOOPK2_else_and_965_nl , LOOPK2_else_and_967_nl , LOOPK2_else_and_969_nl
      , LOOPK2_else_and_971_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1204_nl = ~ LOOPK2_and_61_cse_sva_1;
  assign LOOPK2_if_and_117_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_28_lpi_5, LOOPK2_if_not_1204_nl);
  assign LOOPK2_LOOPK2_nor_29_nl = ~((~(((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_61_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_61_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1009_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1011_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1013_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1015_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1017_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1019_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1021_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1023_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1025_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1027_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1029_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1031_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1033_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1035_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1037_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1039_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1041_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1043_nl = LOOPK2_and_61_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_28_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_28_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_117_nl, {LOOPK2_LOOPK2_nor_29_nl , LOOPK2_else_and_1009_nl ,
      LOOPK2_else_and_1011_nl , LOOPK2_else_and_1013_nl , LOOPK2_else_and_1015_nl
      , LOOPK2_else_and_1017_nl , LOOPK2_else_and_1019_nl , LOOPK2_else_and_1021_nl
      , LOOPK2_else_and_1023_nl , LOOPK2_else_and_1025_nl , LOOPK2_else_and_1027_nl
      , LOOPK2_else_and_1029_nl , LOOPK2_else_and_1031_nl , LOOPK2_else_and_1033_nl
      , LOOPK2_else_and_1035_nl , LOOPK2_else_and_1037_nl , LOOPK2_else_and_1039_nl
      , LOOPK2_else_and_1041_nl , LOOPK2_else_and_1043_nl , operator_38_true_acc_itm_36});
  assign LOOPK2_if_not_1222_nl = ~ LOOPK2_and_60_cse_sva_1;
  assign LOOPK2_if_and_116_nl = MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
      sum_array_27_lpi_5, LOOPK2_if_not_1222_nl);
  assign LOOPK2_LOOPK2_nor_28_nl = ~((~(((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_or_tmp_3)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_or_tmp_2) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_16) | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_130)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_244) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_358) | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_472)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_586) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_700) | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_814)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_928) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_1042) | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_1156)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_1270) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_1384) | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_1498)
      | ((~ LOOPK2_and_60_cse_sva_1) & LOOPK2_else_equal_tmp_1612) | ((~ LOOPK2_and_60_cse_sva_1)
      & LOOPK2_else_equal_tmp_1726) | LOOPK2_else_nor_tmp_1)) | operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_973_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_or_tmp_3
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_975_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_or_tmp_2
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_977_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_16
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_979_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_130
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_981_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_244
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_983_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_358
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_985_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_472
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_987_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_586
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_989_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_700
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_991_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_814
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_993_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_928
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_995_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1042
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_997_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1156
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_999_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1270
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1001_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1384
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1003_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1498
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1005_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1612
      & (~ operator_38_true_acc_itm_36);
  assign LOOPK2_else_and_1007_nl = LOOPK2_and_60_cse_sva_1 & LOOPK2_else_equal_tmp_1726
      & (~ operator_38_true_acc_itm_36);
  assign sum_array_27_lpi_5_dfm_1_mx0w1 = MUX1HOT_v_38_20_2(sum_array_27_sva_2_mx0,
      38'b00000000000000000000000000000000000001, 38'b00000000000000000000000000000000000010,
      38'b00000000000000000000000000000000000011, 38'b00000000000000000000000000000000000100,
      38'b00000000000000000000000000000000000101, 38'b00000000000000000000000000000000000111,
      38'b00000000000000000000000000000000001001, 38'b00000000000000000000000000000000001100,
      38'b00000000000000000000000000000000001111, 38'b00000000000000000000000000000000010100,
      38'b00000000000000000000000000000000011001, 38'b00000000000000000000000000000000100001,
      38'b00000000000000000000000000000000100000, 38'b00000000000000000000000000000000110110,
      38'b00000000000000000000000000000001000110, 38'b00000000000000000000000000000001011010,
      38'b00000000000000000000000000000001110011, 38'b00000000000000000000000000000010010100,
      LOOPK2_if_and_116_nl, {LOOPK2_LOOPK2_nor_28_nl , LOOPK2_else_and_973_nl , LOOPK2_else_and_975_nl
      , LOOPK2_else_and_977_nl , LOOPK2_else_and_979_nl , LOOPK2_else_and_981_nl
      , LOOPK2_else_and_983_nl , LOOPK2_else_and_985_nl , LOOPK2_else_and_987_nl
      , LOOPK2_else_and_989_nl , LOOPK2_else_and_991_nl , LOOPK2_else_and_993_nl
      , LOOPK2_else_and_995_nl , LOOPK2_else_and_997_nl , LOOPK2_else_and_999_nl
      , LOOPK2_else_and_1001_nl , LOOPK2_else_and_1003_nl , LOOPK2_else_and_1005_nl
      , LOOPK2_else_and_1007_nl , operator_38_true_acc_itm_36});
  assign LOOPL1_if_1_unequal_1_itm = ({LOOPK5_k_sva_6 , LOOPK5_k_sva_5_0}) != (z_out_2[6:0]);
  assign LOOPL1_LOOPL1_nor_tmp = ~((z_out_5!=16'b0000000000000000));
  assign LOOPL1_LOOPL1_and_tmp = LOOPK1_endflag_sva & LOOPL1_LOOPL1_nor_tmp;
  assign LOOPK3_if_equal_tmp = LOOPK5_k_sva_5_0 == (z_out_2[6:1]);
  assign LOOPK1_and_stg_3_11_sva_1 = LOOPK1_and_stg_2_3_sva_1 & (cnt_sva[3]);
  assign LOOPK1_and_stg_2_0_sva_1 = LOOPK1_and_stg_1_0_sva_1 & (~ (cnt_sva[2]));
  assign LOOPK1_and_stg_2_1_sva_1 = LOOPK1_and_stg_1_1_sva_1 & (~ (cnt_sva[2]));
  assign LOOPK1_and_stg_2_2_sva_1 = LOOPK1_and_stg_1_2_sva_1 & (~ (cnt_sva[2]));
  assign LOOPK1_and_stg_2_3_sva_1 = LOOPK1_and_stg_1_3_sva_1 & (~ (cnt_sva[2]));
  assign LOOPK1_and_stg_2_4_sva_1 = LOOPK1_and_stg_1_0_sva_1 & (cnt_sva[2]);
  assign LOOPK1_and_stg_2_5_sva_1 = LOOPK1_and_stg_1_1_sva_1 & (cnt_sva[2]);
  assign LOOPK1_and_stg_2_6_sva_1 = LOOPK1_and_stg_1_2_sva_1 & (cnt_sva[2]);
  assign LOOPK1_and_stg_2_7_sva_1 = LOOPK1_and_stg_1_3_sva_1 & (cnt_sva[2]);
  assign LOOPK1_and_stg_1_0_sva_1 = ~((cnt_sva[1:0]!=2'b00));
  assign LOOPK1_and_stg_1_1_sva_1 = (cnt_sva[1:0]==2'b01);
  assign LOOPK1_and_stg_1_2_sva_1 = (cnt_sva[1:0]==2'b10);
  assign LOOPK1_and_stg_1_3_sva_1 = (cnt_sva[1:0]==2'b11);
  assign sum_array_55_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_55_lpi_5,
      or_dcpl_376);
  assign LOOPK2_and_115_cse_sva_1 = LOOPK2_and_stg_4_23_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_0_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_0_lpi_5,
      or_dcpl_374);
  assign LOOPK2_and_114_cse_sva_1 = LOOPK2_and_stg_4_0_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_54_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_54_lpi_5,
      or_dcpl_372);
  assign LOOPK2_and_113_cse_sva_1 = LOOPK2_and_stg_4_22_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_1_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_1_lpi_5,
      or_dcpl_370);
  assign LOOPK2_and_112_cse_sva_1 = LOOPK2_and_stg_4_1_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_53_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_53_lpi_5,
      or_dcpl_368);
  assign LOOPK2_and_111_cse_sva_1 = LOOPK2_and_stg_4_21_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_2_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_2_lpi_5,
      or_dcpl_366);
  assign LOOPK2_and_110_cse_sva_1 = LOOPK2_and_stg_4_2_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_52_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_52_lpi_5,
      or_dcpl_364);
  assign LOOPK2_and_109_cse_sva_1 = LOOPK2_and_stg_4_20_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_3_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_3_lpi_5,
      or_dcpl_362);
  assign LOOPK2_and_108_cse_sva_1 = LOOPK2_and_stg_4_3_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_51_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_51_lpi_5,
      or_dcpl_360);
  assign LOOPK2_and_107_cse_sva_1 = LOOPK2_and_stg_4_19_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_4_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_4_lpi_5,
      or_dcpl_358);
  assign LOOPK2_and_106_cse_sva_1 = LOOPK2_and_stg_4_4_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_50_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_50_lpi_5,
      or_dcpl_356);
  assign LOOPK2_and_105_cse_sva_1 = LOOPK2_and_stg_4_18_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_5_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_5_lpi_5,
      or_dcpl_354);
  assign LOOPK2_and_104_cse_sva_1 = LOOPK2_and_stg_4_5_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_49_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_49_lpi_5,
      or_dcpl_352);
  assign LOOPK2_and_103_cse_sva_1 = LOOPK2_and_stg_4_17_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_6_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_6_lpi_5,
      or_dcpl_350);
  assign LOOPK2_and_102_cse_sva_1 = LOOPK2_and_stg_4_6_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_48_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_48_lpi_5,
      or_dcpl_348);
  assign LOOPK2_and_101_cse_sva_1 = LOOPK2_and_stg_4_16_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_7_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_7_lpi_5,
      or_dcpl_345);
  assign LOOPK2_and_100_cse_sva_1 = LOOPK2_and_stg_4_7_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_47_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_47_lpi_5,
      or_dcpl_342);
  assign LOOPK2_and_99_cse_sva_1 = LOOPK2_and_stg_4_15_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_8_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_8_lpi_5,
      or_dcpl_340);
  assign LOOPK2_and_98_cse_sva_1 = LOOPK2_and_stg_4_8_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_46_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_46_lpi_5,
      or_dcpl_338);
  assign LOOPK2_and_97_cse_sva_1 = LOOPK2_and_stg_4_14_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_9_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_9_lpi_5,
      or_dcpl_336);
  assign LOOPK2_and_96_cse_sva_1 = LOOPK2_and_stg_4_9_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_45_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_45_lpi_5,
      or_dcpl_334);
  assign LOOPK2_and_95_cse_sva_1 = LOOPK2_and_stg_4_13_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_10_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_10_lpi_5,
      or_dcpl_332);
  assign LOOPK2_and_94_cse_sva_1 = LOOPK2_and_stg_4_10_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_44_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_44_lpi_5,
      or_dcpl_330);
  assign LOOPK2_and_93_cse_sva_1 = LOOPK2_and_stg_4_12_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_11_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_11_lpi_5,
      or_dcpl_328);
  assign LOOPK2_and_92_cse_sva_1 = LOOPK2_and_stg_4_11_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_43_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_43_lpi_5,
      or_dcpl_326);
  assign LOOPK2_and_91_cse_sva_1 = LOOPK2_and_stg_4_11_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_12_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_12_lpi_5,
      or_dcpl_323);
  assign LOOPK2_and_90_cse_sva_1 = LOOPK2_and_stg_4_12_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_42_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_42_lpi_5,
      or_dcpl_320);
  assign LOOPK2_and_89_cse_sva_1 = LOOPK2_and_stg_4_10_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_13_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_13_lpi_5,
      or_dcpl_317);
  assign LOOPK2_and_88_cse_sva_1 = LOOPK2_and_stg_4_13_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_41_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_41_lpi_5,
      or_dcpl_314);
  assign LOOPK2_and_87_cse_sva_1 = LOOPK2_and_stg_4_9_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_14_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_14_lpi_5,
      or_dcpl_311);
  assign LOOPK2_and_86_cse_sva_1 = LOOPK2_and_stg_4_14_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_40_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_40_lpi_5,
      or_dcpl_308);
  assign LOOPK2_and_85_cse_sva_1 = LOOPK2_and_stg_4_8_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_15_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_15_lpi_5,
      or_dcpl_304);
  assign LOOPK2_and_84_cse_sva_1 = LOOPK2_and_stg_4_15_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_39_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_39_lpi_5,
      or_dcpl_300);
  assign LOOPK2_and_83_cse_sva_1 = LOOPK2_and_stg_4_7_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_16_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_16_lpi_5,
      or_dcpl_298);
  assign LOOPK2_and_82_cse_sva_1 = LOOPK2_and_stg_4_16_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_38_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_38_lpi_5,
      or_dcpl_296);
  assign LOOPK2_and_81_cse_sva_1 = LOOPK2_and_stg_4_6_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_17_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_17_lpi_5,
      or_dcpl_294);
  assign LOOPK2_and_80_cse_sva_1 = LOOPK2_and_stg_4_17_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_37_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_37_lpi_5,
      or_dcpl_292);
  assign LOOPK2_and_79_cse_sva_1 = LOOPK2_and_stg_4_5_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_18_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_18_lpi_5,
      or_dcpl_289);
  assign LOOPK2_and_78_cse_sva_1 = LOOPK2_and_stg_4_18_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_36_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_36_lpi_5,
      or_dcpl_287);
  assign LOOPK2_and_77_cse_sva_1 = LOOPK2_and_stg_4_4_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_19_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_19_lpi_5,
      or_dcpl_284);
  assign LOOPK2_and_76_cse_sva_1 = LOOPK2_and_stg_4_19_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_35_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_35_lpi_5,
      or_dcpl_282);
  assign LOOPK2_and_75_cse_sva_1 = LOOPK2_and_stg_4_3_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_20_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_20_lpi_5,
      or_dcpl_279);
  assign LOOPK2_and_74_cse_sva_1 = LOOPK2_and_stg_4_20_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_34_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_34_lpi_5,
      or_dcpl_276);
  assign LOOPK2_and_73_cse_sva_1 = LOOPK2_and_stg_4_2_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_21_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_21_lpi_5,
      or_dcpl_272);
  assign LOOPK2_and_72_cse_sva_1 = LOOPK2_and_stg_4_21_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_33_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_33_lpi_5,
      or_dcpl_268);
  assign LOOPK2_and_71_cse_sva_1 = LOOPK2_and_stg_4_1_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_22_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_22_lpi_5,
      or_dcpl_263);
  assign LOOPK2_and_70_cse_sva_1 = LOOPK2_and_stg_4_22_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_32_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_32_lpi_5,
      or_dcpl_260);
  assign LOOPK2_and_69_cse_sva_1 = LOOPK2_and_stg_4_0_sva_1 & (LOOPK5_k_sva_5_0[5]);
  assign sum_array_23_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_23_lpi_5,
      or_dcpl_252);
  assign LOOPK2_and_68_cse_sva_1 = LOOPK2_and_stg_4_23_sva_1 & (~ (LOOPK5_k_sva_5_0[5]));
  assign sum_array_31_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_31_lpi_5,
      or_dcpl_246);
  assign LOOPK2_and_67_cse_sva_1 = LOOPK3_and_stg_3_15_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_24_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_24_lpi_5,
      or_dcpl_243);
  assign LOOPK2_and_66_cse_sva_1 = LOOPK3_and_stg_3_8_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_30_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_30_lpi_5,
      or_dcpl_240);
  assign LOOPK2_and_65_cse_sva_1 = LOOPK3_and_stg_3_14_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_25_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_25_lpi_5,
      or_dcpl_237);
  assign LOOPK2_and_64_cse_sva_1 = LOOPK3_and_stg_3_9_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_29_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_29_lpi_5,
      or_dcpl_234);
  assign LOOPK2_and_63_cse_sva_1 = LOOPK3_and_stg_3_13_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_26_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_26_lpi_5,
      or_dcpl_230);
  assign LOOPK2_and_62_cse_sva_1 = LOOPK3_and_stg_3_10_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_28_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_28_lpi_5,
      or_dcpl_226);
  assign LOOPK2_and_61_cse_sva_1 = LOOPK3_and_stg_3_12_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign sum_array_27_sva_2_mx0 = MUX_v_38_2_2(LOOPK2_acc_ncse_sva_1, sum_array_27_lpi_5,
      or_dcpl_219);
  assign LOOPK2_and_60_cse_sva_1 = LOOPK3_and_stg_3_11_sva_1 & (LOOPK5_k_sva_5_0[5:4]==2'b01);
  assign LOOPK2_else_nor_tmp_1 = ~(LOOPK2_else_LOOPK2_else_and_cse_1 | LOOPK2_else_LOOPK2_else_and_1_cse_1
      | LOOPK2_else_LOOPK2_else_and_2_cse_1 | LOOPK2_else_LOOPK2_else_and_3_cse_1
      | LOOPK2_else_LOOPK2_else_and_4_cse_1 | LOOPK2_else_equal_tmp_16 | LOOPK2_else_equal_tmp_130
      | LOOPK2_else_equal_tmp_244 | LOOPK2_else_equal_tmp_358 | LOOPK2_else_equal_tmp_472
      | LOOPK2_else_equal_tmp_586 | LOOPK2_else_equal_tmp_700 | LOOPK2_else_equal_tmp_814
      | LOOPK2_else_equal_tmp_928 | LOOPK2_else_equal_tmp_1042 | LOOPK2_else_equal_tmp_1156
      | LOOPK2_else_equal_tmp_1270 | LOOPK2_else_equal_tmp_1384 | LOOPK2_else_equal_tmp_1498
      | LOOPK2_else_equal_tmp_1612 | LOOPK2_else_equal_tmp_1726);
  assign LOOPK2_else_equal_tmp_16 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110001);
  assign LOOPK2_else_equal_tmp_130 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110010);
  assign LOOPK2_else_equal_tmp_244 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110011);
  assign LOOPK2_else_equal_tmp_358 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110100);
  assign LOOPK2_else_equal_tmp_472 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110101);
  assign LOOPK2_else_equal_tmp_586 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110110);
  assign LOOPK2_else_equal_tmp_700 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110111);
  assign LOOPK2_else_equal_tmp_814 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111000);
  assign LOOPK2_else_equal_tmp_928 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111001);
  assign LOOPK2_else_equal_tmp_1042 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111010);
  assign LOOPK2_else_equal_tmp_1156 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111011);
  assign LOOPK2_else_equal_tmp_1270 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111100);
  assign LOOPK2_else_equal_tmp_1384 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111101);
  assign LOOPK2_else_equal_tmp_1498 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111110);
  assign LOOPK2_else_equal_tmp_1612 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111111111);
  assign LOOPK2_else_equal_tmp_1726 = ~((LOOPK2_acc_ncse_sva_1!=38'b00000000000000000000000000000000000000));
  assign LOOPK2_else_or_tmp_2 = LOOPK2_else_LOOPK2_else_and_3_cse_1 | LOOPK2_else_LOOPK2_else_and_4_cse_1;
  assign LOOPK2_else_or_tmp_3 = LOOPK2_else_LOOPK2_else_and_cse_1 | LOOPK2_else_LOOPK2_else_and_1_cse_1
      | LOOPK2_else_LOOPK2_else_and_2_cse_1;
  assign LOOPK2_else_LOOPK2_else_and_cse_1 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111101110);
  assign LOOPK2_else_LOOPK2_else_and_1_cse_1 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111101101);
  assign LOOPK2_else_LOOPK2_else_and_2_cse_1 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111101100);
  assign LOOPK2_else_LOOPK2_else_and_3_cse_1 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111110000);
  assign LOOPK2_else_LOOPK2_else_and_4_cse_1 = (LOOPK2_acc_ncse_sva_1==38'b11111111111111111111111111111111101111);
  assign nl_LOOPK2_acc_ncse_sva_1 = LOOPK2_mux_169 - maxn_sva;
  assign LOOPK2_acc_ncse_sva_1 = nl_LOOPK2_acc_ncse_sva_1[37:0];
  assign operator_38_true_operator_38_true_mux_nl = MUX_v_36_56_2((sum_array_0_sva_2_mx0[37:2]),
      (sum_array_1_sva_2_mx0[37:2]), (sum_array_2_sva_2_mx0[37:2]), (sum_array_3_sva_2_mx0[37:2]),
      (sum_array_4_sva_2_mx0[37:2]), (sum_array_5_sva_2_mx0[37:2]), (sum_array_6_sva_2_mx0[37:2]),
      (sum_array_7_sva_2_mx0[37:2]), (sum_array_8_sva_2_mx0[37:2]), (sum_array_9_sva_2_mx0[37:2]),
      (sum_array_10_sva_2_mx0[37:2]), (sum_array_11_sva_2_mx0[37:2]), (sum_array_12_sva_2_mx0[37:2]),
      (sum_array_13_sva_2_mx0[37:2]), (sum_array_14_sva_2_mx0[37:2]), (sum_array_15_sva_2_mx0[37:2]),
      (sum_array_16_sva_2_mx0[37:2]), (sum_array_17_sva_2_mx0[37:2]), (sum_array_18_sva_2_mx0[37:2]),
      (sum_array_19_sva_2_mx0[37:2]), (sum_array_20_sva_2_mx0[37:2]), (sum_array_21_sva_2_mx0[37:2]),
      (sum_array_22_sva_2_mx0[37:2]), (sum_array_23_sva_2_mx0[37:2]), (sum_array_24_sva_2_mx0[37:2]),
      (sum_array_25_sva_2_mx0[37:2]), (sum_array_26_sva_2_mx0[37:2]), (sum_array_27_sva_2_mx0[37:2]),
      (sum_array_28_sva_2_mx0[37:2]), (sum_array_29_sva_2_mx0[37:2]), (sum_array_30_sva_2_mx0[37:2]),
      (sum_array_31_sva_2_mx0[37:2]), (sum_array_32_sva_2_mx0[37:2]), (sum_array_33_sva_2_mx0[37:2]),
      (sum_array_34_sva_2_mx0[37:2]), (sum_array_35_sva_2_mx0[37:2]), (sum_array_36_sva_2_mx0[37:2]),
      (sum_array_37_sva_2_mx0[37:2]), (sum_array_38_sva_2_mx0[37:2]), (sum_array_39_sva_2_mx0[37:2]),
      (sum_array_40_sva_2_mx0[37:2]), (sum_array_41_sva_2_mx0[37:2]), (sum_array_42_sva_2_mx0[37:2]),
      (sum_array_43_sva_2_mx0[37:2]), (sum_array_44_sva_2_mx0[37:2]), (sum_array_45_sva_2_mx0[37:2]),
      (sum_array_46_sva_2_mx0[37:2]), (sum_array_47_sva_2_mx0[37:2]), (sum_array_48_sva_2_mx0[37:2]),
      (sum_array_49_sva_2_mx0[37:2]), (sum_array_50_sva_2_mx0[37:2]), (sum_array_51_sva_2_mx0[37:2]),
      (sum_array_52_sva_2_mx0[37:2]), (sum_array_53_sva_2_mx0[37:2]), (sum_array_54_sva_2_mx0[37:2]),
      (sum_array_55_sva_2_mx0[37:2]), LOOPK5_k_sva_5_0);
  assign nl_operator_38_true_acc_nl = conv_s2u_36_37(operator_38_true_operator_38_true_mux_nl)
      + 37'b0000000000000000000000000000000000101;
  assign operator_38_true_acc_nl = nl_operator_38_true_acc_nl[36:0];
  assign operator_38_true_acc_itm_36 = readslicef_37_1_36(operator_38_true_acc_nl);
  assign LOOPK2_and_stg_4_23_sva_1 = LOOPK3_and_stg_3_7_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_0_sva_1 = LOOPK2_and_stg_3_0_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_22_sva_1 = LOOPK3_and_stg_3_6_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_1_sva_1 = LOOPK3_and_stg_3_1_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_21_sva_1 = LOOPK3_and_stg_3_5_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_2_sva_1 = LOOPK3_and_stg_3_2_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_20_sva_1 = LOOPK3_and_stg_3_4_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_3_sva_1 = LOOPK3_and_stg_3_3_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_19_sva_1 = LOOPK3_and_stg_3_3_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_4_sva_1 = LOOPK3_and_stg_3_4_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_18_sva_1 = LOOPK3_and_stg_3_2_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_5_sva_1 = LOOPK3_and_stg_3_5_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_17_sva_1 = LOOPK3_and_stg_3_1_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_6_sva_1 = LOOPK3_and_stg_3_6_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_16_sva_1 = LOOPK2_and_stg_3_0_sva_1 & (LOOPK5_k_sva_5_0[4]);
  assign LOOPK2_and_stg_4_7_sva_1 = LOOPK3_and_stg_3_7_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_15_sva_1 = LOOPK3_and_stg_3_15_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_8_sva_1 = LOOPK3_and_stg_3_8_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_14_sva_1 = LOOPK3_and_stg_3_14_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_9_sva_1 = LOOPK3_and_stg_3_9_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_13_sva_1 = LOOPK3_and_stg_3_13_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_10_sva_1 = LOOPK3_and_stg_3_10_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_12_sva_1 = LOOPK3_and_stg_3_12_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK2_and_stg_4_11_sva_1 = LOOPK3_and_stg_3_11_sva_1 & (~ (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_and_stg_3_15_sva_1 = LOOPK3_and_stg_2_7_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_8_sva_1 = LOOPK3_and_stg_2_0_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_14_sva_1 = LOOPK3_and_stg_2_6_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_9_sva_1 = LOOPK3_and_stg_2_1_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_13_sva_1 = LOOPK3_and_stg_2_5_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_10_sva_1 = LOOPK3_and_stg_2_2_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_12_sva_1 = LOOPK3_and_stg_2_4_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK3_and_stg_3_11_sva_1 = LOOPK3_and_stg_2_3_sva_1 & (LOOPK5_k_sva_5_0[3]);
  assign LOOPK2_and_stg_3_0_sva_1 = LOOPK3_and_stg_2_0_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_1_sva_1 = LOOPK3_and_stg_2_1_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_2_sva_1 = LOOPK3_and_stg_2_2_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_3_sva_1 = LOOPK3_and_stg_2_3_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_4_sva_1 = LOOPK3_and_stg_2_4_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_5_sva_1 = LOOPK3_and_stg_2_5_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_6_sva_1 = LOOPK3_and_stg_2_6_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_3_7_sva_1 = LOOPK3_and_stg_2_7_sva_1 & (~ (LOOPK5_k_sva_5_0[3]));
  assign LOOPK3_and_stg_2_0_sva_1 = LOOPK3_and_stg_1_0_sva_1 & (~ (LOOPK5_k_sva_5_0[2]));
  assign LOOPK3_and_stg_2_1_sva_1 = LOOPK3_and_stg_1_1_sva_1 & (~ (LOOPK5_k_sva_5_0[2]));
  assign LOOPK3_and_stg_2_2_sva_1 = LOOPK3_and_stg_1_2_sva_1 & (~ (LOOPK5_k_sva_5_0[2]));
  assign LOOPK3_and_stg_2_3_sva_1 = LOOPK3_and_stg_1_3_sva_1 & (~ (LOOPK5_k_sva_5_0[2]));
  assign LOOPK3_and_stg_2_4_sva_1 = LOOPK3_and_stg_1_0_sva_1 & (LOOPK5_k_sva_5_0[2]);
  assign LOOPK3_and_stg_2_5_sva_1 = LOOPK3_and_stg_1_1_sva_1 & (LOOPK5_k_sva_5_0[2]);
  assign LOOPK3_and_stg_2_6_sva_1 = LOOPK3_and_stg_1_2_sva_1 & (LOOPK5_k_sva_5_0[2]);
  assign LOOPK3_and_stg_2_7_sva_1 = LOOPK3_and_stg_1_3_sva_1 & (LOOPK5_k_sva_5_0[2]);
  assign LOOPK3_and_stg_1_0_sva_1 = ~((LOOPK5_k_sva_5_0[1:0]!=2'b00));
  assign LOOPK3_and_stg_1_1_sva_1 = (LOOPK5_k_sva_5_0[1:0]==2'b01);
  assign LOOPK3_and_stg_1_2_sva_1 = (LOOPK5_k_sva_5_0[1:0]==2'b10);
  assign LOOPK3_and_stg_1_3_sva_1 = (LOOPK5_k_sva_5_0[1:0]==2'b11);
  assign LOOPK3_exs_66_0 = ~(LOOPK3_and_stg_3_15_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_68_0 = ~(LOOPK3_and_stg_3_1_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_70_0 = ~(LOOPK3_and_stg_3_14_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_72_0 = ~(LOOPK3_and_stg_3_2_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_74_0 = ~(LOOPK3_and_stg_3_13_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_76_0 = ~(LOOPK3_and_stg_3_3_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_78_0 = ~(LOOPK3_and_stg_3_12_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_80_0 = ~(LOOPK3_and_stg_3_4_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_82_0 = ~(LOOPK3_and_stg_3_11_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_84_0 = ~(LOOPK3_and_stg_3_5_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_86_0 = ~(LOOPK3_and_stg_3_10_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_88_0 = ~(LOOPK3_and_stg_3_6_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_90_0 = ~(LOOPK3_and_stg_3_9_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_92_0 = ~(LOOPK3_and_stg_3_7_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_94_0 = ~(LOOPK3_and_stg_3_8_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_96_0 = ~(LOOPK3_and_stg_3_8_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_98_0 = ~(LOOPK3_and_stg_3_7_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_100_0 = ~(LOOPK3_and_stg_3_9_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_102_0 = ~(LOOPK3_and_stg_3_6_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_104_0 = ~(LOOPK3_and_stg_3_10_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_106_0 = ~(LOOPK3_and_stg_3_5_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_108_0 = ~(LOOPK3_and_stg_3_11_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_110_0 = ~(LOOPK3_and_stg_3_4_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_112_0 = ~(LOOPK3_and_stg_3_12_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_114_0 = ~(LOOPK3_and_stg_3_3_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_116_0 = ~(LOOPK3_and_stg_3_13_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_118_0 = ~(LOOPK3_and_stg_3_2_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_120_0 = ~(LOOPK3_and_stg_3_14_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_122_0 = ~(LOOPK3_and_stg_3_1_sva_1 & (LOOPK5_k_sva_5_0[4]));
  assign LOOPK3_exs_124_0 = ~(LOOPK3_and_stg_3_15_sva_1 & (~ (LOOPK5_k_sva_5_0[4])));
  assign LOOPK3_exs_126_0 = ~(LOOPK3_and_stg_2_0_sva_1 & (LOOPK5_k_sva_5_0[4:3]==2'b10));
  assign nl_operator_4_false_acc_psp_sva_1 = conv_u2s_4_5(head) + 5'b11111;
  assign operator_4_false_acc_psp_sva_1 = nl_operator_4_false_acc_psp_sva_1[4:0];
  assign LOOPK2_mux_169 = MUX_v_38_56_2(sum_array_0_lpi_5, sum_array_1_lpi_5, sum_array_2_lpi_5,
      sum_array_3_lpi_5, sum_array_4_lpi_5, sum_array_5_lpi_5, sum_array_6_lpi_5,
      sum_array_7_lpi_5, sum_array_8_lpi_5, sum_array_9_lpi_5, sum_array_10_lpi_5,
      sum_array_11_lpi_5, sum_array_12_lpi_5, sum_array_13_lpi_5, sum_array_14_lpi_5,
      sum_array_15_lpi_5, sum_array_16_lpi_5, sum_array_17_lpi_5, sum_array_18_lpi_5,
      sum_array_19_lpi_5, sum_array_20_lpi_5, sum_array_21_lpi_5, sum_array_22_lpi_5,
      sum_array_23_lpi_5, sum_array_24_lpi_5, sum_array_25_lpi_5, sum_array_26_lpi_5,
      sum_array_27_lpi_5, sum_array_28_lpi_5, sum_array_29_lpi_5, sum_array_30_lpi_5,
      sum_array_31_lpi_5, sum_array_32_lpi_5, sum_array_33_lpi_5, sum_array_34_lpi_5,
      sum_array_35_lpi_5, sum_array_36_lpi_5, sum_array_37_lpi_5, sum_array_38_lpi_5,
      sum_array_39_lpi_5, sum_array_40_lpi_5, sum_array_41_lpi_5, sum_array_42_lpi_5,
      sum_array_43_lpi_5, sum_array_44_lpi_5, sum_array_45_lpi_5, sum_array_46_lpi_5,
      sum_array_47_lpi_5, sum_array_48_lpi_5, sum_array_49_lpi_5, sum_array_50_lpi_5,
      sum_array_51_lpi_5, sum_array_52_lpi_5, sum_array_53_lpi_5, sum_array_54_lpi_5,
      sum_array_55_lpi_5, LOOPK5_k_sva_5_0);
  assign LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp = ~((LOOPI1_i_sva != (operator_4_false_acc_psp_sva_1[3:0]))
      | (operator_4_false_acc_psp_sva_1[4]));
  assign LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp = ~((LOOPJ1_j_sva != (z_out_2[5:0]))
      | (z_out_2[6]));
  assign LOOPK2_if_1_equal_1_tmp = LOOPK5_k_sva_5_0 == (z_out_1[5:0]);
  assign LOOPK4_LOOPK4_if_1_and_tmp = LOOPK2_if_1_equal_1_tmp & (z_out_1[8:6]==3'b000);
  assign LOOPK3_if_unequal_tmp = LOOPK5_k_sva_5_0 != (z_out_2[6:1]);
  assign and_363_cse = (~ LOOPK4_LOOPK4_if_1_and_tmp) & (fsm_output[11]);
  assign and_dcpl_83 = (~ (LOOPK5_k_sva_5_0[5])) & (LOOPK5_k_sva_5_0[0]);
  assign and_dcpl_84 = and_dcpl_83 & (~ (LOOPK5_k_sva_5_0[2]));
  assign and_dcpl_85 = (LOOPK5_k_sva_5_0[1]) & (LOOPK5_k_sva_5_0[3]);
  assign and_dcpl_86 = and_dcpl_85 & (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_215 = (LOOPK5_k_sva_5_0[5]) | (~ (LOOPK5_k_sva_5_0[0]));
  assign or_dcpl_216 = or_dcpl_215 | (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_217 = ~((LOOPK5_k_sva_5_0[1]) & (LOOPK5_k_sva_5_0[3]));
  assign or_dcpl_218 = or_dcpl_217 | (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_219 = or_dcpl_218 | or_dcpl_216;
  assign and_dcpl_90 = ~((LOOPK5_k_sva_5_0[5]) | (LOOPK5_k_sva_5_0[0]));
  assign and_dcpl_91 = and_dcpl_90 & (LOOPK5_k_sva_5_0[2]);
  assign and_dcpl_92 = (~ (LOOPK5_k_sva_5_0[1])) & (LOOPK5_k_sva_5_0[3]);
  assign and_dcpl_93 = and_dcpl_92 & (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_222 = (LOOPK5_k_sva_5_0[5]) | (LOOPK5_k_sva_5_0[0]);
  assign or_dcpl_223 = or_dcpl_222 | (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_224 = (LOOPK5_k_sva_5_0[1]) | (~ (LOOPK5_k_sva_5_0[3]));
  assign or_dcpl_225 = or_dcpl_224 | (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_226 = or_dcpl_225 | or_dcpl_223;
  assign and_dcpl_97 = and_dcpl_90 & (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_229 = or_dcpl_222 | (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_230 = or_dcpl_218 | or_dcpl_229;
  assign and_dcpl_101 = and_dcpl_83 & (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_233 = or_dcpl_215 | (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_234 = or_dcpl_225 | or_dcpl_233;
  assign or_dcpl_237 = or_dcpl_225 | or_dcpl_216;
  assign or_dcpl_240 = or_dcpl_218 | or_dcpl_223;
  assign or_dcpl_243 = or_dcpl_225 | or_dcpl_229;
  assign or_dcpl_246 = or_dcpl_218 | or_dcpl_233;
  assign or_dcpl_247 = (~ LOOPK1_slc_cnt_5_0_10_itm) | LOOPK1_slc_cnt_5_0_66_itm;
  assign or_dcpl_248 = (~ LOOPK1_and_stg_2_7_sva) | LOOPK1_slc_cnt_5_0_9_itm;
  assign and_dcpl_115 = LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm);
  assign and_dcpl_116 = LOOPK1_and_stg_2_7_sva & (~ LOOPK1_slc_cnt_5_0_9_itm);
  assign and_dcpl_118 = (LOOPK5_k_sva_5_0[1]) & (~ (LOOPK5_k_sva_5_0[3]));
  assign and_dcpl_119 = and_dcpl_118 & (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_250 = (~ (LOOPK5_k_sva_5_0[1])) | (LOOPK5_k_sva_5_0[3]);
  assign or_dcpl_251 = or_dcpl_250 | (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_252 = or_dcpl_251 | or_dcpl_233;
  assign or_dcpl_253 = LOOPK1_slc_cnt_5_0_10_itm | (~ LOOPK1_slc_cnt_5_0_66_itm);
  assign or_dcpl_254 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_0_sva);
  assign and_dcpl_121 = (~ LOOPK1_slc_cnt_5_0_10_itm) & LOOPK1_slc_cnt_5_0_66_itm;
  assign and_dcpl_122 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_0_sva;
  assign and_dcpl_124 = (LOOPK5_k_sva_5_0[5]) & (~ (LOOPK5_k_sva_5_0[0]));
  assign and_dcpl_125 = and_dcpl_124 & (~ (LOOPK5_k_sva_5_0[2]));
  assign and_dcpl_126 = ~((LOOPK5_k_sva_5_0[1]) | (LOOPK5_k_sva_5_0[3]));
  assign and_dcpl_127 = and_dcpl_126 & (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_256 = (~ (LOOPK5_k_sva_5_0[5])) | (LOOPK5_k_sva_5_0[0]);
  assign or_dcpl_257 = or_dcpl_256 | (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_258 = (LOOPK5_k_sva_5_0[1]) | (LOOPK5_k_sva_5_0[3]);
  assign or_dcpl_259 = or_dcpl_258 | (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_260 = or_dcpl_259 | or_dcpl_257;
  assign or_dcpl_261 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_6_sva);
  assign and_dcpl_129 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_6_sva;
  assign or_dcpl_263 = or_dcpl_251 | or_dcpl_223;
  assign or_dcpl_264 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_1_sva);
  assign and_dcpl_132 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_1_sva;
  assign and_dcpl_134 = (LOOPK5_k_sva_5_0[5]) & (LOOPK5_k_sva_5_0[0]);
  assign and_dcpl_135 = and_dcpl_134 & (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_266 = ~((LOOPK5_k_sva_5_0[5]) & (LOOPK5_k_sva_5_0[0]));
  assign or_dcpl_267 = or_dcpl_266 | (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_268 = or_dcpl_259 | or_dcpl_267;
  assign or_dcpl_269 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_5_sva);
  assign and_dcpl_137 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_5_sva;
  assign and_dcpl_139 = and_dcpl_126 & (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_271 = or_dcpl_258 | (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_272 = or_dcpl_271 | or_dcpl_233;
  assign or_dcpl_273 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_2_sva);
  assign and_dcpl_141 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_2_sva;
  assign and_dcpl_143 = and_dcpl_118 & (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_275 = or_dcpl_250 | (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_276 = or_dcpl_275 | or_dcpl_257;
  assign or_dcpl_277 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_4_sva);
  assign and_dcpl_145 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_4_sva;
  assign or_dcpl_279 = or_dcpl_271 | or_dcpl_223;
  assign or_dcpl_280 = LOOPK1_slc_cnt_5_0_9_itm | (~ LOOPK1_and_stg_2_3_sva);
  assign and_dcpl_148 = (~ LOOPK1_slc_cnt_5_0_9_itm) & LOOPK1_and_stg_2_3_sva;
  assign or_dcpl_282 = or_dcpl_275 | or_dcpl_267;
  assign or_dcpl_284 = or_dcpl_251 | or_dcpl_216;
  assign and_dcpl_154 = and_dcpl_124 & (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_286 = or_dcpl_256 | (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_287 = or_dcpl_259 | or_dcpl_286;
  assign or_dcpl_289 = or_dcpl_251 | or_dcpl_229;
  assign and_dcpl_159 = and_dcpl_134 & (LOOPK5_k_sva_5_0[2]);
  assign or_dcpl_291 = or_dcpl_266 | (~ (LOOPK5_k_sva_5_0[2]));
  assign or_dcpl_292 = or_dcpl_259 | or_dcpl_291;
  assign or_dcpl_294 = or_dcpl_271 | or_dcpl_216;
  assign or_dcpl_296 = or_dcpl_275 | or_dcpl_286;
  assign or_dcpl_298 = or_dcpl_271 | or_dcpl_229;
  assign or_dcpl_300 = or_dcpl_275 | or_dcpl_291;
  assign or_dcpl_301 = (~ LOOPK1_and_stg_3_15_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_169 = LOOPK1_and_stg_3_15_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign and_dcpl_171 = and_dcpl_85 & (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_303 = or_dcpl_217 | (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_304 = or_dcpl_303 | or_dcpl_233;
  assign or_dcpl_305 = (~ LOOPK1_and_stg_3_8_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_173 = LOOPK1_and_stg_3_8_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign and_dcpl_175 = and_dcpl_92 & (~ (LOOPK5_k_sva_5_0[4]));
  assign or_dcpl_307 = or_dcpl_224 | (LOOPK5_k_sva_5_0[4]);
  assign or_dcpl_308 = or_dcpl_307 | or_dcpl_257;
  assign or_dcpl_309 = (~ LOOPK1_and_stg_3_14_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_177 = LOOPK1_and_stg_3_14_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_311 = or_dcpl_303 | or_dcpl_223;
  assign or_dcpl_312 = (~ LOOPK1_and_stg_3_9_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_180 = LOOPK1_and_stg_3_9_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_314 = or_dcpl_307 | or_dcpl_267;
  assign or_dcpl_315 = (~ LOOPK1_and_stg_3_13_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_183 = LOOPK1_and_stg_3_13_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_317 = or_dcpl_307 | or_dcpl_233;
  assign or_dcpl_318 = (~ LOOPK1_and_stg_3_10_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_186 = LOOPK1_and_stg_3_10_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_320 = or_dcpl_303 | or_dcpl_257;
  assign or_dcpl_321 = (~ LOOPK1_and_stg_3_12_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_189 = LOOPK1_and_stg_3_12_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_323 = or_dcpl_307 | or_dcpl_223;
  assign or_dcpl_324 = (~ LOOPK1_and_stg_3_11_sva) | LOOPK1_slc_cnt_5_0_10_itm;
  assign and_dcpl_192 = LOOPK1_and_stg_3_11_sva & (~ LOOPK1_slc_cnt_5_0_10_itm);
  assign or_dcpl_326 = or_dcpl_303 | or_dcpl_267;
  assign or_dcpl_328 = or_dcpl_303 | or_dcpl_216;
  assign or_dcpl_330 = or_dcpl_307 | or_dcpl_286;
  assign or_dcpl_332 = or_dcpl_303 | or_dcpl_229;
  assign or_dcpl_334 = or_dcpl_307 | or_dcpl_291;
  assign or_dcpl_336 = or_dcpl_307 | or_dcpl_216;
  assign or_dcpl_338 = or_dcpl_303 | or_dcpl_286;
  assign or_dcpl_340 = or_dcpl_307 | or_dcpl_229;
  assign or_dcpl_342 = or_dcpl_303 | or_dcpl_291;
  assign or_dcpl_343 = LOOPK1_slc_cnt_5_0_10_itm | LOOPK1_slc_cnt_5_0_66_itm;
  assign and_dcpl_211 = ~(LOOPK1_slc_cnt_5_0_10_itm | LOOPK1_slc_cnt_5_0_66_itm);
  assign or_dcpl_345 = or_dcpl_275 | or_dcpl_233;
  assign or_dcpl_346 = ~(LOOPK1_slc_cnt_5_0_10_itm & LOOPK1_slc_cnt_5_0_66_itm);
  assign and_dcpl_214 = LOOPK1_slc_cnt_5_0_10_itm & LOOPK1_slc_cnt_5_0_66_itm;
  assign or_dcpl_348 = or_dcpl_271 | or_dcpl_257;
  assign or_dcpl_350 = or_dcpl_275 | or_dcpl_223;
  assign or_dcpl_352 = or_dcpl_271 | or_dcpl_267;
  assign or_dcpl_354 = or_dcpl_259 | or_dcpl_233;
  assign or_dcpl_356 = or_dcpl_251 | or_dcpl_257;
  assign or_dcpl_358 = or_dcpl_259 | or_dcpl_223;
  assign or_dcpl_360 = or_dcpl_251 | or_dcpl_267;
  assign or_dcpl_362 = or_dcpl_275 | or_dcpl_216;
  assign or_dcpl_364 = or_dcpl_271 | or_dcpl_286;
  assign or_dcpl_366 = or_dcpl_275 | or_dcpl_229;
  assign or_dcpl_368 = or_dcpl_271 | or_dcpl_291;
  assign or_dcpl_370 = or_dcpl_259 | or_dcpl_216;
  assign or_dcpl_372 = or_dcpl_251 | or_dcpl_286;
  assign or_dcpl_374 = or_dcpl_259 | or_dcpl_229;
  assign or_dcpl_376 = or_dcpl_251 | or_dcpl_291;
  assign and_dcpl_245 = ~((LOOPL2_l_sva[4:3]!=2'b00));
  assign and_dcpl_246 = and_dcpl_245 & (LOOPL2_l_sva[5]);
  assign and_dcpl_247 = ~((LOOPL2_l_sva[1:0]!=2'b00));
  assign and_dcpl_248 = and_dcpl_247 & (~ (LOOPL2_l_sva[2]));
  assign and_dcpl_251 = (LOOPL2_l_sva[4:3]==2'b11);
  assign and_dcpl_252 = and_dcpl_251 & (~ (LOOPL2_l_sva[5]));
  assign and_dcpl_253 = (LOOPL2_l_sva[1:0]==2'b10);
  assign and_dcpl_254 = and_dcpl_253 & (LOOPL2_l_sva[2]);
  assign and_dcpl_256 = and_dcpl_253 & (~ (LOOPL2_l_sva[2]));
  assign and_dcpl_258 = and_dcpl_247 & (LOOPL2_l_sva[2]);
  assign and_dcpl_264 = (LOOPL2_l_sva[4:3]==2'b01);
  assign and_dcpl_265 = and_dcpl_264 & (LOOPL2_l_sva[5]);
  assign and_dcpl_267 = (LOOPL2_l_sva[4:3]==2'b10);
  assign and_dcpl_268 = and_dcpl_267 & (~ (LOOPL2_l_sva[5]));
  assign and_dcpl_276 = and_dcpl_267 & (LOOPL2_l_sva[5]);
  assign and_dcpl_278 = and_dcpl_264 & (~ (LOOPL2_l_sva[5]));
  assign and_dcpl_286 = and_dcpl_251 & (LOOPL2_l_sva[5]);
  assign and_dcpl_288 = and_dcpl_245 & (~ (LOOPL2_l_sva[5]));
  assign and_dcpl_295 = (LOOPL2_l_sva[1:0]==2'b11);
  assign and_dcpl_296 = and_dcpl_295 & (LOOPL2_l_sva[2]);
  assign and_dcpl_300 = (LOOPL2_l_sva[1:0]==2'b01);
  assign and_dcpl_301 = and_dcpl_300 & (~ (LOOPL2_l_sva[2]));
  assign and_dcpl_303 = and_dcpl_300 & (LOOPL2_l_sva[2]);
  assign and_dcpl_305 = and_dcpl_295 & (~ (LOOPL2_l_sva[2]));
  assign and_dcpl_348 = ~((fsm_output[11:10]!=2'b00));
  assign and_671_cse = (fsm_output[9:4]==6'b000000);
  assign or_tmp_553 = (fsm_output[2]) | (fsm_output[11]);
  assign LOOPK5_mux_cse = MUX_v_6_2_2(LOOPK5_k_sva_5_0, (LOOPL2_l_sva[5:0]), fsm_output[10]);
  assign or_tmp_759 = (LOOPL2_l_sva[4:0]!=5'b00000) | nand_58_cse;
  assign or_tmp_766 = (LOOPL2_l_sva[4:0]!=5'b00010) | nand_58_cse;
  assign or_tmp_773 = (LOOPL2_l_sva[4:0]!=5'b00100) | nand_58_cse;
  assign or_tmp_780 = (LOOPL2_l_sva[4:0]!=5'b00110) | nand_58_cse;
  assign or_tmp_787 = (LOOPL2_l_sva[4:0]!=5'b01000) | nand_58_cse;
  assign or_tmp_794 = (LOOPL2_l_sva[4:0]!=5'b01010) | nand_58_cse;
  assign or_tmp_801 = (LOOPL2_l_sva[4:0]!=5'b01100) | nand_58_cse;
  assign or_tmp_808 = (LOOPL2_l_sva[4:0]!=5'b01110) | nand_58_cse;
  assign or_tmp_815 = (LOOPL2_l_sva[3:0]!=4'b0000) | nand_75_cse;
  assign or_tmp_822 = (LOOPL2_l_sva[3:0]!=4'b0010) | nand_75_cse;
  assign or_tmp_829 = (LOOPL2_l_sva[3:0]!=4'b0100) | nand_75_cse;
  assign or_tmp_836 = (LOOPL2_l_sva[3:0]!=4'b0110) | nand_75_cse;
  assign or_tmp_843 = (LOOPL2_l_sva[2:0]!=3'b000) | nand_84_cse;
  assign or_tmp_850 = (LOOPL2_l_sva[2:0]!=3'b010) | nand_84_cse;
  assign or_tmp_857 = (LOOPL2_l_sva[1:0]!=2'b00) | nand_55_cse;
  assign or_tmp_868 = nand_22_cse | nor_14_cse;
  assign nand_108_cse = ~((LOOPK5_k_sva_5_0[4]) & or_1735_cse);
  assign or_tmp_873 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0000) | nand_108_cse;
  assign or_tmp_878 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01110) | nor_14_cse;
  assign or_tmp_883 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0001) | nand_108_cse;
  assign or_tmp_888 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01101) | nor_14_cse;
  assign or_tmp_893 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0010) | nand_108_cse;
  assign or_tmp_898 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01100) | nor_14_cse;
  assign or_tmp_903 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0011) | nand_108_cse;
  assign or_tmp_908 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01011) | nor_14_cse;
  assign or_tmp_913 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0100) | nand_108_cse;
  assign or_tmp_918 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01010) | nor_14_cse;
  assign or_tmp_923 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0101) | nand_108_cse;
  assign or_tmp_928 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01001) | nor_14_cse;
  assign or_tmp_933 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0110) | nand_108_cse;
  assign or_tmp_938 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01000) | nor_14_cse;
  assign or_tmp_943 = nand_31_cse | nand_108_cse;
  assign or_tmp_948 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00111) | nor_14_cse;
  assign nand_117_cse = ~((LOOPK5_k_sva_5_0[4:3]==2'b11) & or_1735_cse);
  assign or_tmp_953 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b000) | nand_117_cse;
  assign or_tmp_958 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00110) | nor_14_cse;
  assign or_tmp_963 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b001) | nand_117_cse;
  assign or_tmp_968 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00101) | nor_14_cse;
  assign or_tmp_973 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b010) | nand_117_cse;
  assign or_tmp_978 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00100) | nor_14_cse;
  assign or_tmp_983 = nand_44_cse | nand_117_cse;
  assign or_tmp_988 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00011) | nor_14_cse;
  assign nand_122_cse = ~((LOOPK5_k_sva_5_0[4:2]==3'b111) & or_1735_cse);
  assign or_tmp_993 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[1:0]!=2'b00) | nand_122_cse;
  assign or_tmp_998 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00010) | nor_14_cse;
  assign or_tmp_1003 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[1:0]!=2'b01) | nand_122_cse;
  assign or_tmp_1008 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00001) |
      nor_14_cse;
  assign or_tmp_1012 = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[0]) | (~((LOOPK5_k_sva_5_0[4:1]==4'b1111)
      & or_1735_cse));
  assign not_tmp_714 = ~((fsm_output[10:9]!=2'b00));
  assign or_1731_nl = (z_out_2[7]) | LOOPL1_if_1_unequal_1_itm | not_tmp_714;
  assign mux_tmp_46 = MUX_s_1_2_2(not_tmp_714, or_1731_nl, fsm_output[3]);
  assign or_1253_itm = (((z_out_2[7]) | LOOPL1_if_1_unequal_1_itm) & (fsm_output[3]))
      | (fsm_output[12]);
  assign LOOPL1_mux_1_itm = MUX_v_16_64_2((q_channel_data_sva[15:0]), (q_channel_data_sva[31:16]),
      (q_channel_data_sva[47:32]), (q_channel_data_sva[63:48]), (q_channel_data_sva[79:64]),
      (q_channel_data_sva[95:80]), (q_channel_data_sva[111:96]), (q_channel_data_sva[127:112]),
      (q_channel_data_sva[143:128]), (q_channel_data_sva[159:144]), (q_channel_data_sva[175:160]),
      (q_channel_data_sva[191:176]), (q_channel_data_sva[207:192]), (q_channel_data_sva[223:208]),
      (q_channel_data_sva[239:224]), (q_channel_data_sva[255:240]), (q_channel_data_sva[271:256]),
      (q_channel_data_sva[287:272]), (q_channel_data_sva[303:288]), (q_channel_data_sva[319:304]),
      (q_channel_data_sva[335:320]), (q_channel_data_sva[351:336]), (q_channel_data_sva[367:352]),
      (q_channel_data_sva[383:368]), (q_channel_data_sva[399:384]), (q_channel_data_sva[415:400]),
      (q_channel_data_sva[431:416]), (q_channel_data_sva[447:432]), (q_channel_data_sva[463:448]),
      (q_channel_data_sva[479:464]), (q_channel_data_sva[495:480]), (q_channel_data_sva[511:496]),
      (q_channel_data_sva[527:512]), (q_channel_data_sva[543:528]), (q_channel_data_sva[559:544]),
      (q_channel_data_sva[575:560]), (q_channel_data_sva[591:576]), (q_channel_data_sva[607:592]),
      (q_channel_data_sva[623:608]), (q_channel_data_sva[639:624]), (q_channel_data_sva[655:640]),
      (q_channel_data_sva[671:656]), (q_channel_data_sva[687:672]), (q_channel_data_sva[703:688]),
      (q_channel_data_sva[719:704]), (q_channel_data_sva[735:720]), (q_channel_data_sva[751:736]),
      (q_channel_data_sva[767:752]), (q_channel_data_sva[783:768]), (q_channel_data_sva[799:784]),
      (q_channel_data_sva[815:800]), (q_channel_data_sva[831:816]), (q_channel_data_sva[847:832]),
      (q_channel_data_sva[863:848]), (q_channel_data_sva[879:864]), (q_channel_data_sva[895:880]),
      (q_channel_data_sva[911:896]), (q_channel_data_sva[927:912]), (q_channel_data_sva[943:928]),
      (q_channel_data_sva[959:944]), (q_channel_data_sva[975:960]), (q_channel_data_sva[991:976]),
      (q_channel_data_sva[1007:992]), (q_channel_data_sva[1023:1008]), LOOPK5_k_sva_5_0);
  always @(posedge clk) begin
    if ( run_wen & LOOPI1_i_or_cse ) begin
      LOOPI1_i_sva <= MUX_v_4_2_2(4'b0000, operator_4_false_acc_nl, LOOPI1_i_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & ((fsm_output[14]) | LOOPI1_i_or_cse) ) begin
      LOOPJ1_j_sva <= MUX_v_6_2_2(6'b000000, z_out, not_254_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[12]) ) begin
      dout_chan_rsci_idat <= z_out_4;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((~ LOOPK1_and_60_itm) & (fsm_output[4])))) )
        begin
      sum_array_27_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_27_lpi_5, {and_675_nl , and_677_nl , and_679_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_12_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_28_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_28_lpi_5, {and_684_nl , and_686_nl , and_688_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_10_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_26_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_26_lpi_5, {and_693_nl , and_695_nl , and_697_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_13_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_29_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_29_lpi_5, {and_702_nl , and_704_nl , and_706_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_9_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_25_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_25_lpi_5, {and_711_nl , and_713_nl , and_715_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_14_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_30_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_30_lpi_5, {and_720_nl , and_722_nl , and_724_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_8_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_24_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_24_lpi_5, {and_729_nl , and_731_nl , and_733_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | (((~(LOOPK1_and_stg_3_15_sva & LOOPK1_slc_cnt_5_0_10_itm))
        | LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4])))) ) begin
      sum_array_31_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_31_lpi_5, {and_738_nl , and_740_nl , and_742_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_248 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_23_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_23_lpi_5, {and_747_nl , and_749_nl , and_751_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_254 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_32_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_32_lpi_5, {and_756_nl , and_758_nl , and_760_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_261 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_22_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_22_lpi_5, {and_765_nl , and_767_nl , and_769_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_264 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_33_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_33_lpi_5, {and_774_nl , and_776_nl , and_778_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_269 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_21_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_21_lpi_5, {and_783_nl , and_785_nl , and_787_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_273 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_34_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_34_lpi_5, {and_792_nl , and_794_nl , and_796_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_277 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_20_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_20_lpi_5, {and_801_nl , and_803_nl , and_805_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_280 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_35_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_35_lpi_5, {and_810_nl , and_812_nl , and_814_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_280 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_19_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_19_lpi_5, {and_819_nl , and_821_nl , and_823_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_277 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_36_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_36_lpi_5, {and_828_nl , and_830_nl , and_832_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_273 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_18_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_18_lpi_5, {and_837_nl , and_839_nl , and_841_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_269 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_37_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_37_lpi_5, {and_846_nl , and_848_nl , and_850_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_264 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_17_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_17_lpi_5, {and_855_nl , and_857_nl , and_859_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_261 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_38_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_38_lpi_5, {and_864_nl , and_866_nl , and_868_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_254 | or_dcpl_247) & (fsm_output[4]))))
        ) begin
      sum_array_16_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_16_lpi_5, {and_873_nl , and_875_nl , and_877_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_248 | or_dcpl_253) & (fsm_output[4]))))
        ) begin
      sum_array_39_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_39_lpi_5, {and_882_nl , and_884_nl , and_886_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_301 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_15_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_15_lpi_5, {and_891_nl , and_893_nl , and_895_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_305 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_40_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_40_lpi_5, {and_900_nl , and_902_nl , and_904_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_309 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_14_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_14_lpi_5, {and_909_nl , and_911_nl , and_913_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_312 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_41_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_41_lpi_5, {and_918_nl , and_920_nl , and_922_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_315 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_13_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_13_lpi_5, {and_927_nl , and_929_nl , and_931_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_318 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_42_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_42_lpi_5, {and_936_nl , and_938_nl , and_940_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_321 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_12_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_12_lpi_5, {and_945_nl , and_947_nl , and_949_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_324 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_43_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_43_lpi_5, {and_954_nl , and_956_nl , and_958_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_324 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_11_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_11_lpi_5, {and_963_nl , and_965_nl , and_967_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_321 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_44_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_44_lpi_5, {and_972_nl , and_974_nl , and_976_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_318 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_10_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_10_lpi_5, {and_981_nl , and_983_nl , and_985_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_315 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_45_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_45_lpi_5, {and_990_nl , and_992_nl , and_994_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_312 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_9_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_9_lpi_5, {and_999_nl , and_1001_nl , and_1003_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_309 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_46_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_46_lpi_5, {and_1008_nl , and_1010_nl , and_1012_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_305 | LOOPK1_slc_cnt_5_0_66_itm) &
        (fsm_output[4])))) ) begin
      sum_array_8_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_8_lpi_5, {and_1017_nl , and_1019_nl , and_1021_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_301 | (~ LOOPK1_slc_cnt_5_0_66_itm))
        & (fsm_output[4])))) ) begin
      sum_array_47_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_47_lpi_5, {and_1026_nl , and_1028_nl , and_1030_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_248 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_7_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_7_lpi_5, {and_1035_nl , and_1037_nl , and_1039_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_254 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_48_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_48_lpi_5, {and_1044_nl , and_1046_nl , and_1048_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_261 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_6_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_6_lpi_5, {and_1053_nl , and_1055_nl , and_1057_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_264 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_49_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_49_lpi_5, {and_1062_nl , and_1064_nl , and_1066_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_269 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_5_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_5_lpi_5, {and_1071_nl , and_1073_nl , and_1075_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_273 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_50_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_50_lpi_5, {and_1080_nl , and_1082_nl , and_1084_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_277 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_4_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_4_lpi_5, {and_1089_nl , and_1091_nl , and_1093_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_280 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_51_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_51_lpi_5, {and_1098_nl , and_1100_nl , and_1102_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_280 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_3_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_3_lpi_5, {and_1107_nl , and_1109_nl , and_1111_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_277 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_52_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_52_lpi_5, {and_1116_nl , and_1118_nl , and_1120_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_273 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_2_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_2_lpi_5, {and_1125_nl , and_1127_nl , and_1129_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_269 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_53_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_53_lpi_5, {and_1134_nl , and_1136_nl , and_1138_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_264 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_1_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_1_lpi_5, {and_1143_nl , and_1145_nl , and_1147_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_261 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_54_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_54_lpi_5, {and_1152_nl , and_1154_nl , and_1156_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_254 | or_dcpl_343) & (fsm_output[4]))))
        ) begin
      sum_array_0_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_0_lpi_5, {and_1161_nl , and_1163_nl , and_1165_nl});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(and_671_cse | ((or_dcpl_248 | or_dcpl_346) & (fsm_output[4]))))
        ) begin
      sum_array_55_lpi_3 <= MUX1HOT_v_38_3_2((signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          z_out_6, sum_array_55_lpi_5, {and_1170_nl , and_1172_nl , and_1174_nl});
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_nl) & run_wen ) begin
      data_out_32_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_60_nl, z_out_3, and_1178_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(nand_22_cse & (~((LOOPL2_l_sva[5:0]==6'b011110) & (fsm_output[10])))))
        & run_wen ) begin
      data_out_30_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_61_nl, z_out_3, and_1185_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_6_nl) & run_wen ) begin
      data_out_34_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_62_nl, z_out_3, and_1192_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01110)) & ((LOOPL2_l_sva[5:0]!=6'b011100)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_28_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_63_nl, z_out_3, and_1199_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_7_nl) & run_wen ) begin
      data_out_36_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_64_nl, z_out_3, and_1206_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01101)) & ((LOOPL2_l_sva[5:0]!=6'b011010)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_26_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_65_nl, z_out_3, and_1213_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_8_nl) & run_wen ) begin
      data_out_38_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_66_nl, z_out_3, and_1220_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01100)) & ((LOOPL2_l_sva[5:0]!=6'b011000)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_24_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_67_nl, z_out_3, and_1227_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_9_nl) & run_wen ) begin
      data_out_40_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_68_nl, z_out_3, and_1234_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01011)) & ((LOOPL2_l_sva[5:0]!=6'b010110)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_22_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_69_nl, z_out_3, and_1241_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_10_nl) & run_wen ) begin
      data_out_42_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_70_nl, z_out_3, and_1248_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01010)) & ((LOOPL2_l_sva[5:0]!=6'b010100)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_20_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_71_nl, z_out_3, and_1255_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_11_nl) & run_wen ) begin
      data_out_44_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_72_nl, z_out_3, and_1262_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01001)) & ((LOOPL2_l_sva[5:0]!=6'b010010)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_18_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_73_nl, z_out_3, and_1269_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_12_nl) & run_wen ) begin
      data_out_46_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_74_nl, z_out_3, and_1276_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b01000)) & ((LOOPL2_l_sva[5:0]!=6'b010000)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_16_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_75_nl, z_out_3, and_1283_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_13_nl) & run_wen ) begin
      data_out_48_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_76_nl, z_out_3, and_1290_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00111)) & ((LOOPL2_l_sva[5:0]!=6'b001110)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_14_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_77_nl, z_out_3, and_1297_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_14_nl) & run_wen ) begin
      data_out_50_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_78_nl, z_out_3, and_1304_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00110)) & ((LOOPL2_l_sva[5:0]!=6'b001100)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_12_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_79_nl, z_out_3, and_1311_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_15_nl) & run_wen ) begin
      data_out_52_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_80_nl, z_out_3, and_1318_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00101)) & ((LOOPL2_l_sva[5:0]!=6'b001010)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_10_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_81_nl, z_out_3, and_1325_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_16_nl) & run_wen ) begin
      data_out_54_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_82_nl, z_out_3, and_1332_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00100)) & ((LOOPL2_l_sva[5:0]!=6'b001000)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_8_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_83_nl, z_out_3, and_1339_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_17_nl) & run_wen ) begin
      data_out_56_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_84_nl, z_out_3, and_1346_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00011)) & ((LOOPL2_l_sva[5:0]!=6'b000110)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_6_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_85_nl, z_out_3, and_1353_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_18_nl) & run_wen ) begin
      data_out_58_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_86_nl, z_out_3, and_1360_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00010)) & ((LOOPL2_l_sva[5:0]!=6'b000100)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_4_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_87_nl, z_out_3, and_1367_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_19_nl) & run_wen ) begin
      data_out_60_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_88_nl, z_out_3, and_1374_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~(((~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[4:0]!=5'b00001)) & ((LOOPL2_l_sva[5:0]!=6'b000010)
        | (~ (fsm_output[10]))))) & run_wen ) begin
      data_out_2_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_89_nl, z_out_3, and_1381_nl);
    end
  end
  always @(posedge clk) begin
    if ( (((fsm_output[7]) & (LOOPK5_k_sva_5_0[4:0]==5'b11111)) | (~((LOOPL2_l_sva[1:0]!=2'b10)
        | nand_55_cse))) & run_wen ) begin
      data_out_62_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_90_nl, z_out_3, and_1388_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_20_nl) & run_wen ) begin
      data_out_31_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_152_nl, z_out_3, and_1395_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_21_nl) & run_wen ) begin
      data_out_33_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_153_nl, z_out_3, and_1402_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_22_nl) & run_wen ) begin
      data_out_29_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_154_nl, z_out_3, and_1409_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_23_nl) & run_wen ) begin
      data_out_35_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_155_nl, z_out_3, and_1416_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_24_nl) & run_wen ) begin
      data_out_27_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_156_nl, z_out_3, and_1423_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_25_nl) & run_wen ) begin
      data_out_37_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_157_nl, z_out_3, and_1430_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_26_nl) & run_wen ) begin
      data_out_25_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_158_nl, z_out_3, and_1437_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_27_nl) & run_wen ) begin
      data_out_39_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_159_nl, z_out_3, and_1444_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_28_nl) & run_wen ) begin
      data_out_23_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_160_nl, z_out_3, and_1451_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_29_nl) & run_wen ) begin
      data_out_41_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_161_nl, z_out_3, and_1458_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_30_nl) & run_wen ) begin
      data_out_21_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_162_nl, z_out_3, and_1465_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_31_nl) & run_wen ) begin
      data_out_43_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_163_nl, z_out_3, and_1472_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_32_nl) & run_wen ) begin
      data_out_19_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_164_nl, z_out_3, and_1479_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_33_nl) & run_wen ) begin
      data_out_45_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_165_nl, z_out_3, and_1486_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_34_nl) & run_wen ) begin
      data_out_17_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_166_nl, z_out_3, and_1493_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_35_nl) & run_wen ) begin
      data_out_47_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_167_nl, z_out_3, and_1500_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_36_nl) & run_wen ) begin
      data_out_15_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_168_nl, z_out_3, and_1507_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_37_nl) & run_wen ) begin
      data_out_49_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_169_nl, z_out_3, and_1514_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_38_nl) & run_wen ) begin
      data_out_13_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_170_nl, z_out_3, and_1521_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_39_nl) & run_wen ) begin
      data_out_51_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_171_nl, z_out_3, and_1528_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_40_nl) & run_wen ) begin
      data_out_11_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_172_nl, z_out_3, and_1535_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_41_nl) & run_wen ) begin
      data_out_53_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_173_nl, z_out_3, and_1542_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_42_nl) & run_wen ) begin
      data_out_9_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_174_nl, z_out_3, and_1549_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_43_nl) & run_wen ) begin
      data_out_55_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_175_nl, z_out_3, and_1556_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_44_nl) & run_wen ) begin
      data_out_7_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_176_nl, z_out_3, and_1563_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_45_nl) & run_wen ) begin
      data_out_57_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_177_nl, z_out_3, and_1570_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_46_nl) & run_wen ) begin
      data_out_5_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_178_nl, z_out_3, and_1577_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_47_nl) & run_wen ) begin
      data_out_59_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_179_nl, z_out_3, and_1584_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_48_nl) & run_wen ) begin
      data_out_3_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_180_nl, z_out_3, and_1591_nl);
    end
  end
  always @(posedge clk) begin
    if ( (~ mux_49_nl) & run_wen ) begin
      data_out_61_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_181_nl, z_out_3, and_1598_nl);
    end
  end
  always @(posedge clk) begin
    if ( ((~(((LOOPL2_l_sva[3:0]!=4'b0001) | (~ (fsm_output[10])) | (LOOPL2_l_sva[5:4]!=2'b00))
        & (~(or_1735_cse & (fsm_output[7]))))) | and_2155_cse) & run_wen & (~((nor_14_cse
        & (fsm_output[7])) | ((~ LOOPK1_endflag_sva) & (fsm_output[8])))) ) begin
      data_out_1_lpi_3 <= ~(MUX_v_16_2_2(nor_402_nl, 16'b1111111111111111, or_1744_nl));
    end
  end
  always @(posedge clk) begin
    if ( (((LOOPL2_l_sva[5:0]==6'b111111) & (fsm_output[10])) | ((fsm_output[7])
        & (LOOPK5_k_sva_5_0[4:0]==5'b11111) & or_1735_cse)) & run_wen ) begin
      data_out_63_lpi_3 <= MUX_v_16_2_2(LOOPK3_and_183_nl, z_out_3, and_1614_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_q_chan2_rsci_oswt_cse <= 1'b0;
      reg_k_chan2_rsci_oswt_cse <= 1'b0;
      reg_v_chan2_rsci_oswt_cse <= 1'b0;
      reg_dout_chan_rsci_oswt_cse <= 1'b0;
      LOOPK1_endflag_sva <= 1'b0;
      LOOPK5_k_sva_6 <= 1'b0;
      LOOPL2_l_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( rst ) begin
      reg_q_chan2_rsci_oswt_cse <= 1'b0;
      reg_k_chan2_rsci_oswt_cse <= 1'b0;
      reg_v_chan2_rsci_oswt_cse <= 1'b0;
      reg_dout_chan_rsci_oswt_cse <= 1'b0;
      LOOPK1_endflag_sva <= 1'b0;
      LOOPK5_k_sva_6 <= 1'b0;
      LOOPL2_l_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( run_wen ) begin
      reg_q_chan2_rsci_oswt_cse <= ~((LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp & (fsm_output[15]))
          | (~((fsm_output[14]) | (fsm_output[0]) | (fsm_output[15]))) | (LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp
          & (fsm_output[14])));
      reg_k_chan2_rsci_oswt_cse <= (fsm_output[1]) | (fsm_output[4]);
      reg_v_chan2_rsci_oswt_cse <= and_363_cse | (fsm_output[8]);
      reg_dout_chan_rsci_oswt_cse <= fsm_output[12];
      LOOPK1_endflag_sva <= LOOPK1_endflag_mux1h_2_nl | (~((fsm_output[12]) | (fsm_output[3])
          | (fsm_output[7])));
      LOOPK5_k_sva_6 <= LOOPL1_l_LOOPL1_l_mux_nl & LOOPK5_k_nor_seb;
      LOOPL2_l_sva <= MUX_v_32_2_2(32'b00000000000000000000000000000000, LOOPL2_acc_1_nl,
          (fsm_output[10]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      cnt_sva <= 8'b00000000;
    end
    else if ( rst ) begin
      cnt_sva <= 8'b00000000;
    end
    else if ( ((((z_out_5!=16'b0000000000000000) | (~ LOOPK1_endflag_sva)) & nor_169_cse
        & (fsm_output[3])) | (fsm_output[15]) | (fsm_output[0]) | (fsm_output[1])
        | (fsm_output[13]) | (fsm_output[14]) | (fsm_output[16]) | (fsm_output[12]))
        & run_wen ) begin
      cnt_sva <= MUX_v_8_2_2(8'b00000000, (z_out_1[7:0]), cnt_nor_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (((fsm_output[5:2]==4'b0000)) | and_1639_rgt) ) begin
      maxn_sva <= MUX_v_38_2_2(38'b10000000000000000000000000000000000000, (signext_38_13(LOOPL1_ac_int_cctor_sva[37:25])),
          and_1639_rgt);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[4:2]==3'b000) ) begin
      q_channel_data_sva <= q_chan2_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b110111)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_55_lpi_5 <= MUX_v_38_2_2(sum_array_55_lpi_5_dfm_1_mx0w1, sum_array_55_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_177_cse & nor_178_cse) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_0_lpi_5 <= MUX_v_38_2_2(sum_array_0_lpi_5_dfm_1_mx0w1, sum_array_0_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b110110)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_54_lpi_5 <= MUX_v_38_2_2(sum_array_54_lpi_5_dfm_1_mx0w1, sum_array_54_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (~ (LOOPK5_k_sva_5_0[3]))
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_1_lpi_5 <= MUX_v_38_2_2(sum_array_1_lpi_5_dfm_1_mx0w1, sum_array_1_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_53_lpi_5 <= MUX_v_38_2_2(sum_array_53_lpi_5_dfm_1_mx0w1, sum_array_53_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_177_cse & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_2_lpi_5 <= MUX_v_38_2_2(sum_array_2_lpi_5_dfm_1_mx0w1, sum_array_2_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_52_lpi_5 <= MUX_v_38_2_2(sum_array_52_lpi_5_dfm_1_mx0w1, sum_array_52_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b0011) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_3_lpi_5 <= MUX_v_38_2_2(sum_array_3_lpi_5_dfm_1_mx0w1, sum_array_3_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b110011)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_51_lpi_5 <= MUX_v_38_2_2(sum_array_51_lpi_5_dfm_1_mx0w1, sum_array_51_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_4_lpi_5 <= MUX_v_38_2_2(sum_array_4_lpi_5_dfm_1_mx0w1, sum_array_4_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b11))
        | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_50_lpi_5 <= MUX_v_38_2_2(sum_array_50_lpi_5_dfm_1_mx0w1, sum_array_50_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_5_lpi_5 <= MUX_v_38_2_2(sum_array_5_lpi_5_dfm_1_mx0w1, sum_array_5_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_49_lpi_5 <= MUX_v_38_2_2(sum_array_49_lpi_5_dfm_1_mx0w1, sum_array_49_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b0110) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_6_lpi_5 <= MUX_v_38_2_2(sum_array_6_lpi_5_dfm_1_mx0w1, sum_array_6_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b11)) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_48_lpi_5 <= MUX_v_38_2_2(sum_array_48_lpi_5_dfm_1_mx0w1, sum_array_48_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b0111) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_7_lpi_5 <= MUX_v_38_2_2(sum_array_7_lpi_5_dfm_1_mx0w1, sum_array_7_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b101111)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_47_lpi_5 <= MUX_v_38_2_2(sum_array_47_lpi_5_dfm_1_mx0w1, sum_array_47_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_240_cse & (LOOPK5_k_sva_5_0[3]) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_8_lpi_5 <= MUX_v_38_2_2(sum_array_8_lpi_5_dfm_1_mx0w1, sum_array_8_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b101110)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_46_lpi_5 <= MUX_v_38_2_2(sum_array_46_lpi_5_dfm_1_mx0w1, sum_array_46_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (LOOPK5_k_sva_5_0[3])
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_9_lpi_5 <= MUX_v_38_2_2(sum_array_9_lpi_5_dfm_1_mx0w1, sum_array_9_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_45_lpi_5 <= MUX_v_38_2_2(sum_array_45_lpi_5_dfm_1_mx0w1, sum_array_45_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_240_cse & (LOOPK5_k_sva_5_0[3])
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_10_lpi_5 <= MUX_v_38_2_2(sum_array_10_lpi_5_dfm_1_mx0w1, sum_array_10_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_44_lpi_5 <= MUX_v_38_2_2(sum_array_44_lpi_5_dfm_1_mx0w1, sum_array_44_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b1011) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_11_lpi_5 <= MUX_v_38_2_2(sum_array_11_lpi_5_dfm_1_mx0w1, sum_array_11_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b101011)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_43_lpi_5 <= MUX_v_38_2_2(sum_array_43_lpi_5_dfm_1_mx0w1, sum_array_43_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_12_lpi_5 <= MUX_v_38_2_2(sum_array_12_lpi_5_dfm_1_mx0w1, sum_array_12_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_240_cse & (LOOPK5_k_sva_5_0[5:3]==3'b101))
        | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_42_lpi_5 <= MUX_v_38_2_2(sum_array_42_lpi_5_dfm_1_mx0w1, sum_array_42_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & nor_178_cse) | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_13_lpi_5 <= MUX_v_38_2_2(sum_array_13_lpi_5_dfm_1_mx0w1, sum_array_13_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_41_lpi_5 <= MUX_v_38_2_2(sum_array_41_lpi_5_dfm_1_mx0w1, sum_array_41_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b1110) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_14_lpi_5 <= MUX_v_38_2_2(sum_array_14_lpi_5_dfm_1_mx0w1, sum_array_14_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_240_cse & (LOOPK5_k_sva_5_0[5:3]==3'b101)) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_40_lpi_5 <= MUX_v_38_2_2(sum_array_40_lpi_5_dfm_1_mx0w1, sum_array_40_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[3:0]==4'b1111) & nor_178_cse) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_15_lpi_5 <= MUX_v_38_2_2(sum_array_15_lpi_5_dfm_1_mx0w1, sum_array_15_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b100111)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_39_lpi_5 <= MUX_v_38_2_2(sum_array_39_lpi_5_dfm_1_mx0w1, sum_array_39_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b01)) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_16_lpi_5 <= MUX_v_38_2_2(sum_array_16_lpi_5_dfm_1_mx0w1, sum_array_16_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b100110)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_38_lpi_5 <= MUX_v_38_2_2(sum_array_38_lpi_5_dfm_1_mx0w1, sum_array_38_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (~ (LOOPK5_k_sva_5_0[5]))) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_17_lpi_5 <= MUX_v_38_2_2(sum_array_17_lpi_5_dfm_1_mx0w1, sum_array_17_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_37_lpi_5 <= MUX_v_38_2_2(sum_array_37_lpi_5_dfm_1_mx0w1, sum_array_37_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b01))
        | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_18_lpi_5 <= MUX_v_38_2_2(sum_array_18_lpi_5_dfm_1_mx0w1, sum_array_18_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_36_lpi_5 <= MUX_v_38_2_2(sum_array_36_lpi_5_dfm_1_mx0w1, sum_array_36_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b010011)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_19_lpi_5 <= MUX_v_38_2_2(sum_array_19_lpi_5_dfm_1_mx0w1, sum_array_19_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b100011)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_35_lpi_5 <= MUX_v_38_2_2(sum_array_35_lpi_5_dfm_1_mx0w1, sum_array_35_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (~ (LOOPK5_k_sva_5_0[5]))) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_20_lpi_5 <= MUX_v_38_2_2(sum_array_20_lpi_5_dfm_1_mx0w1, sum_array_20_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b10))
        | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_34_lpi_5 <= MUX_v_38_2_2(sum_array_34_lpi_5_dfm_1_mx0w1, sum_array_34_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (~ (LOOPK5_k_sva_5_0[3]))
        & (LOOPK5_k_sva_5_0[4]) & (~ (LOOPK5_k_sva_5_0[5]))) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_21_lpi_5 <= MUX_v_38_2_2(sum_array_21_lpi_5_dfm_1_mx0w1, sum_array_21_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (~ (LOOPK5_k_sva_5_0[3]))
        & (~ (LOOPK5_k_sva_5_0[4])) & (LOOPK5_k_sva_5_0[5])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_33_lpi_5 <= MUX_v_38_2_2(sum_array_33_lpi_5_dfm_1_mx0w1, sum_array_33_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b010110)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_22_lpi_5 <= MUX_v_38_2_2(sum_array_22_lpi_5_dfm_1_mx0w1, sum_array_22_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_177_cse & (LOOPK5_k_sva_5_0[5:4]==2'b10)) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_32_lpi_5 <= MUX_v_38_2_2(sum_array_32_lpi_5_dfm_1_mx0w1, sum_array_32_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b010111)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_23_lpi_5 <= MUX_v_38_2_2(sum_array_23_lpi_5_dfm_1_mx0w1, sum_array_23_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b011111)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_31_lpi_5 <= MUX_v_38_2_2(sum_array_31_lpi_5_dfm_1_mx0w1, sum_array_31_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & nor_240_cse & (LOOPK5_k_sva_5_0[5:3]==3'b011)) | (fsm_output[11])
        | (fsm_output[2])) & run_wen ) begin
      sum_array_24_lpi_5 <= MUX_v_38_2_2(sum_array_24_lpi_5_dfm_1_mx0w1, sum_array_24_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b011110)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_30_lpi_5 <= MUX_v_38_2_2(sum_array_30_lpi_5_dfm_1_mx0w1, sum_array_30_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (~ (LOOPK5_k_sva_5_0[2])) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[5])) & (LOOPK5_k_sva_5_0[4])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_25_lpi_5 <= MUX_v_38_2_2(sum_array_25_lpi_5_dfm_1_mx0w1, sum_array_25_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (LOOPK5_k_sva_5_0[0]) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[5])) & (LOOPK5_k_sva_5_0[4])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_29_lpi_5 <= MUX_v_38_2_2(sum_array_29_lpi_5_dfm_1_mx0w1, sum_array_29_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0[1]) & nor_240_cse & (LOOPK5_k_sva_5_0[5:3]==3'b011))
        | (fsm_output[11]) | (fsm_output[2])) & run_wen ) begin
      sum_array_26_lpi_5 <= MUX_v_38_2_2(sum_array_26_lpi_5_dfm_1_mx0w1, sum_array_26_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((nor_174_cse & (~ (LOOPK5_k_sva_5_0[0])) & (LOOPK5_k_sva_5_0[2]) & (LOOPK5_k_sva_5_0[3])
        & (~ (LOOPK5_k_sva_5_0[5])) & (LOOPK5_k_sva_5_0[4])) | (fsm_output[11]) |
        (fsm_output[2])) & run_wen ) begin
      sum_array_28_lpi_5 <= MUX_v_38_2_2(sum_array_28_lpi_5_dfm_1_mx0w1, sum_array_28_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( ((and_2169_cse & (LOOPK5_k_sva_5_0==6'b011011)) | (fsm_output[11]) | (fsm_output[2]))
        & run_wen ) begin
      sum_array_27_lpi_5 <= MUX_v_38_2_2(sum_array_27_lpi_5_dfm_1_mx0w1, sum_array_27_lpi_3,
          or_tmp_553);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~((fsm_output[3]) | (fsm_output[10]))) ) begin
      k_channel_data_sva <= MUX_v_1024_2_2(k_chan2_rsci_idat_mxwt, v_chan2_rsci_idat_mxwt,
          fsm_output[9]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPK5_k_sva_5_0 <= 6'b000000;
    end
    else if ( rst ) begin
      LOOPK5_k_sva_5_0 <= 6'b000000;
    end
    else if ( (mux_52_nl | (fsm_output[4]) | (fsm_output[15]) | (fsm_output[1]) |
        (fsm_output[14]) | (fsm_output[2]) | (fsm_output[16]) | (fsm_output[0]) |
        (fsm_output[12])) & run_wen ) begin
      LOOPK5_k_sva_5_0 <= MUX_v_6_2_2(6'b000000, LOOPL1_l_LOOPL1_l_mux_1_nl, and_2822_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen ) begin
      LOOPL1_ac_int_cctor_sva <= MUX_v_38_2_2(38'b00000000000000000000000000000000000000,
          LOOPL1_acc_nl, (fsm_output[3]));
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[11:7]==5'b00000) ) begin
      LOOPJ1_sum2_1_sva <= MUX_v_16_2_2(16'b0000000000000000, LOOPJ1_sum2_mux_nl,
          not_370_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPK1_slc_cnt_5_0_66_itm <= 1'b0;
      LOOPK1_and_stg_3_15_sva <= 1'b0;
      LOOPK1_slc_cnt_5_0_10_itm <= 1'b0;
      LOOPK1_and_stg_3_14_sva <= 1'b0;
      LOOPK1_and_stg_3_13_sva <= 1'b0;
      LOOPK1_and_stg_3_12_sva <= 1'b0;
      LOOPK1_and_60_itm <= 1'b0;
      LOOPK1_and_stg_3_10_sva <= 1'b0;
      LOOPK1_and_stg_3_9_sva <= 1'b0;
      LOOPK1_and_stg_3_8_sva <= 1'b0;
      LOOPK1_and_stg_3_11_sva <= 1'b0;
      LOOPK1_and_stg_2_0_sva <= 1'b0;
      LOOPK1_slc_cnt_5_0_9_itm <= 1'b0;
      LOOPK1_and_stg_2_1_sva <= 1'b0;
      LOOPK1_and_stg_2_2_sva <= 1'b0;
      LOOPK1_and_stg_2_3_sva <= 1'b0;
      LOOPK1_and_stg_2_4_sva <= 1'b0;
      LOOPK1_and_stg_2_5_sva <= 1'b0;
      LOOPK1_and_stg_2_6_sva <= 1'b0;
      LOOPK1_and_stg_2_7_sva <= 1'b0;
    end
    else if ( rst ) begin
      LOOPK1_slc_cnt_5_0_66_itm <= 1'b0;
      LOOPK1_and_stg_3_15_sva <= 1'b0;
      LOOPK1_slc_cnt_5_0_10_itm <= 1'b0;
      LOOPK1_and_stg_3_14_sva <= 1'b0;
      LOOPK1_and_stg_3_13_sva <= 1'b0;
      LOOPK1_and_stg_3_12_sva <= 1'b0;
      LOOPK1_and_60_itm <= 1'b0;
      LOOPK1_and_stg_3_10_sva <= 1'b0;
      LOOPK1_and_stg_3_9_sva <= 1'b0;
      LOOPK1_and_stg_3_8_sva <= 1'b0;
      LOOPK1_and_stg_3_11_sva <= 1'b0;
      LOOPK1_and_stg_2_0_sva <= 1'b0;
      LOOPK1_slc_cnt_5_0_9_itm <= 1'b0;
      LOOPK1_and_stg_2_1_sva <= 1'b0;
      LOOPK1_and_stg_2_2_sva <= 1'b0;
      LOOPK1_and_stg_2_3_sva <= 1'b0;
      LOOPK1_and_stg_2_4_sva <= 1'b0;
      LOOPK1_and_stg_2_5_sva <= 1'b0;
      LOOPK1_and_stg_2_6_sva <= 1'b0;
      LOOPK1_and_stg_2_7_sva <= 1'b0;
    end
    else if ( LOOPK1_and_61_cse ) begin
      LOOPK1_slc_cnt_5_0_66_itm <= cnt_sva[5];
      LOOPK1_and_stg_3_15_sva <= LOOPK1_and_stg_2_7_sva_1 & (cnt_sva[3]);
      LOOPK1_slc_cnt_5_0_10_itm <= cnt_sva[4];
      LOOPK1_and_stg_3_14_sva <= LOOPK1_and_stg_2_6_sva_1 & (cnt_sva[3]);
      LOOPK1_and_stg_3_13_sva <= LOOPK1_and_stg_2_5_sva_1 & (cnt_sva[3]);
      LOOPK1_and_stg_3_12_sva <= LOOPK1_and_stg_2_4_sva_1 & (cnt_sva[3]);
      LOOPK1_and_60_itm <= LOOPK1_and_stg_3_11_sva_1 & (cnt_sva[5:4]==2'b01);
      LOOPK1_and_stg_3_10_sva <= LOOPK1_and_stg_2_2_sva_1 & (cnt_sva[3]);
      LOOPK1_and_stg_3_9_sva <= LOOPK1_and_stg_2_1_sva_1 & (cnt_sva[3]);
      LOOPK1_and_stg_3_8_sva <= LOOPK1_and_stg_2_0_sva_1 & (cnt_sva[3]);
      LOOPK1_and_stg_3_11_sva <= LOOPK1_and_stg_3_11_sva_1;
      LOOPK1_and_stg_2_0_sva <= LOOPK1_and_stg_2_0_sva_1;
      LOOPK1_slc_cnt_5_0_9_itm <= cnt_sva[3];
      LOOPK1_and_stg_2_1_sva <= LOOPK1_and_stg_2_1_sva_1;
      LOOPK1_and_stg_2_2_sva <= LOOPK1_and_stg_2_2_sva_1;
      LOOPK1_and_stg_2_3_sva <= LOOPK1_and_stg_2_3_sva_1;
      LOOPK1_and_stg_2_4_sva <= LOOPK1_and_stg_2_4_sva_1;
      LOOPK1_and_stg_2_5_sva <= LOOPK1_and_stg_2_5_sva_1;
      LOOPK1_and_stg_2_6_sva <= LOOPK1_and_stg_2_6_sva_1;
      LOOPK1_and_stg_2_7_sva <= LOOPK1_and_stg_2_7_sva_1;
    end
  end
  always @(posedge clk) begin
    if ( (~((~((LOOPL2_l_sva[5:0]==6'b000000))) & (fsm_output[10]))) & (~((fsm_output[11])
        | (fsm_output[9]) | (fsm_output[12]))) & (~ (fsm_output[13])) & run_wen )
        begin
      data_out_0_lpi_6 <= MUX_v_16_2_2(16'b0000000000000000, z_out_3, data_out_nand_nl);
    end
  end
  assign nl_operator_4_false_acc_nl = LOOPI1_i_sva + 4'b0001;
  assign operator_4_false_acc_nl = nl_operator_4_false_acc_nl[3:0];
  assign LOOPI1_i_not_1_nl = ~ (fsm_output[0]);
  assign not_254_nl = ~ LOOPI1_i_or_cse;
  assign and_675_nl = LOOPK1_and_60_itm & (fsm_output[4]);
  assign and_677_nl = and_dcpl_86 & and_dcpl_84 & (fsm_output[9]);
  assign and_679_nl = or_dcpl_219 & (fsm_output[9]);
  assign and_684_nl = LOOPK1_and_stg_3_12_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_686_nl = and_dcpl_93 & and_dcpl_91 & (fsm_output[9]);
  assign and_688_nl = or_dcpl_226 & (fsm_output[9]);
  assign and_693_nl = LOOPK1_and_stg_3_10_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_695_nl = and_dcpl_86 & and_dcpl_97 & (fsm_output[9]);
  assign and_697_nl = or_dcpl_230 & (fsm_output[9]);
  assign and_702_nl = LOOPK1_and_stg_3_13_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_704_nl = and_dcpl_93 & and_dcpl_101 & (fsm_output[9]);
  assign and_706_nl = or_dcpl_234 & (fsm_output[9]);
  assign and_711_nl = LOOPK1_and_stg_3_9_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_713_nl = and_dcpl_93 & and_dcpl_84 & (fsm_output[9]);
  assign and_715_nl = or_dcpl_237 & (fsm_output[9]);
  assign and_720_nl = LOOPK1_and_stg_3_14_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_722_nl = and_dcpl_86 & and_dcpl_91 & (fsm_output[9]);
  assign and_724_nl = or_dcpl_240 & (fsm_output[9]);
  assign and_729_nl = LOOPK1_and_stg_3_8_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_731_nl = and_dcpl_93 & and_dcpl_97 & (fsm_output[9]);
  assign and_733_nl = or_dcpl_243 & (fsm_output[9]);
  assign and_738_nl = LOOPK1_and_stg_3_15_sva & LOOPK1_slc_cnt_5_0_10_itm & (~ LOOPK1_slc_cnt_5_0_66_itm)
      & (fsm_output[4]);
  assign and_740_nl = and_dcpl_86 & and_dcpl_101 & (fsm_output[9]);
  assign and_742_nl = or_dcpl_246 & (fsm_output[9]);
  assign and_747_nl = and_dcpl_116 & and_dcpl_115 & (fsm_output[4]);
  assign and_749_nl = and_dcpl_119 & and_dcpl_101 & (fsm_output[9]);
  assign and_751_nl = or_dcpl_252 & (fsm_output[9]);
  assign and_756_nl = and_dcpl_122 & and_dcpl_121 & (fsm_output[4]);
  assign and_758_nl = and_dcpl_127 & and_dcpl_125 & (fsm_output[9]);
  assign and_760_nl = or_dcpl_260 & (fsm_output[9]);
  assign and_765_nl = and_dcpl_129 & and_dcpl_115 & (fsm_output[4]);
  assign and_767_nl = and_dcpl_119 & and_dcpl_91 & (fsm_output[9]);
  assign and_769_nl = or_dcpl_263 & (fsm_output[9]);
  assign and_774_nl = and_dcpl_132 & and_dcpl_121 & (fsm_output[4]);
  assign and_776_nl = and_dcpl_127 & and_dcpl_135 & (fsm_output[9]);
  assign and_778_nl = or_dcpl_268 & (fsm_output[9]);
  assign and_783_nl = and_dcpl_137 & and_dcpl_115 & (fsm_output[4]);
  assign and_785_nl = and_dcpl_139 & and_dcpl_101 & (fsm_output[9]);
  assign and_787_nl = or_dcpl_272 & (fsm_output[9]);
  assign and_792_nl = and_dcpl_141 & and_dcpl_121 & (fsm_output[4]);
  assign and_794_nl = and_dcpl_143 & and_dcpl_125 & (fsm_output[9]);
  assign and_796_nl = or_dcpl_276 & (fsm_output[9]);
  assign and_801_nl = and_dcpl_145 & and_dcpl_115 & (fsm_output[4]);
  assign and_803_nl = and_dcpl_139 & and_dcpl_91 & (fsm_output[9]);
  assign and_805_nl = or_dcpl_279 & (fsm_output[9]);
  assign and_810_nl = and_dcpl_148 & and_dcpl_121 & (fsm_output[4]);
  assign and_812_nl = and_dcpl_143 & and_dcpl_135 & (fsm_output[9]);
  assign and_814_nl = or_dcpl_282 & (fsm_output[9]);
  assign and_819_nl = and_dcpl_148 & and_dcpl_115 & (fsm_output[4]);
  assign and_821_nl = and_dcpl_119 & and_dcpl_84 & (fsm_output[9]);
  assign and_823_nl = or_dcpl_284 & (fsm_output[9]);
  assign and_828_nl = and_dcpl_145 & and_dcpl_121 & (fsm_output[4]);
  assign and_830_nl = and_dcpl_127 & and_dcpl_154 & (fsm_output[9]);
  assign and_832_nl = or_dcpl_287 & (fsm_output[9]);
  assign and_837_nl = and_dcpl_141 & and_dcpl_115 & (fsm_output[4]);
  assign and_839_nl = and_dcpl_119 & and_dcpl_97 & (fsm_output[9]);
  assign and_841_nl = or_dcpl_289 & (fsm_output[9]);
  assign and_846_nl = and_dcpl_137 & and_dcpl_121 & (fsm_output[4]);
  assign and_848_nl = and_dcpl_127 & and_dcpl_159 & (fsm_output[9]);
  assign and_850_nl = or_dcpl_292 & (fsm_output[9]);
  assign and_855_nl = and_dcpl_132 & and_dcpl_115 & (fsm_output[4]);
  assign and_857_nl = and_dcpl_139 & and_dcpl_84 & (fsm_output[9]);
  assign and_859_nl = or_dcpl_294 & (fsm_output[9]);
  assign and_864_nl = and_dcpl_129 & and_dcpl_121 & (fsm_output[4]);
  assign and_866_nl = and_dcpl_143 & and_dcpl_154 & (fsm_output[9]);
  assign and_868_nl = or_dcpl_296 & (fsm_output[9]);
  assign and_873_nl = and_dcpl_122 & and_dcpl_115 & (fsm_output[4]);
  assign and_875_nl = and_dcpl_139 & and_dcpl_97 & (fsm_output[9]);
  assign and_877_nl = or_dcpl_298 & (fsm_output[9]);
  assign and_882_nl = and_dcpl_116 & and_dcpl_121 & (fsm_output[4]);
  assign and_884_nl = and_dcpl_143 & and_dcpl_159 & (fsm_output[9]);
  assign and_886_nl = or_dcpl_300 & (fsm_output[9]);
  assign and_891_nl = and_dcpl_169 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_893_nl = and_dcpl_171 & and_dcpl_101 & (fsm_output[9]);
  assign and_895_nl = or_dcpl_304 & (fsm_output[9]);
  assign and_900_nl = and_dcpl_173 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_902_nl = and_dcpl_175 & and_dcpl_125 & (fsm_output[9]);
  assign and_904_nl = or_dcpl_308 & (fsm_output[9]);
  assign and_909_nl = and_dcpl_177 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_911_nl = and_dcpl_171 & and_dcpl_91 & (fsm_output[9]);
  assign and_913_nl = or_dcpl_311 & (fsm_output[9]);
  assign and_918_nl = and_dcpl_180 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_920_nl = and_dcpl_175 & and_dcpl_135 & (fsm_output[9]);
  assign and_922_nl = or_dcpl_314 & (fsm_output[9]);
  assign and_927_nl = and_dcpl_183 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_929_nl = and_dcpl_175 & and_dcpl_101 & (fsm_output[9]);
  assign and_931_nl = or_dcpl_317 & (fsm_output[9]);
  assign and_936_nl = and_dcpl_186 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_938_nl = and_dcpl_171 & and_dcpl_125 & (fsm_output[9]);
  assign and_940_nl = or_dcpl_320 & (fsm_output[9]);
  assign and_945_nl = and_dcpl_189 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_947_nl = and_dcpl_175 & and_dcpl_91 & (fsm_output[9]);
  assign and_949_nl = or_dcpl_323 & (fsm_output[9]);
  assign and_954_nl = and_dcpl_192 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_956_nl = and_dcpl_171 & and_dcpl_135 & (fsm_output[9]);
  assign and_958_nl = or_dcpl_326 & (fsm_output[9]);
  assign and_963_nl = and_dcpl_192 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_965_nl = and_dcpl_171 & and_dcpl_84 & (fsm_output[9]);
  assign and_967_nl = or_dcpl_328 & (fsm_output[9]);
  assign and_972_nl = and_dcpl_189 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_974_nl = and_dcpl_175 & and_dcpl_154 & (fsm_output[9]);
  assign and_976_nl = or_dcpl_330 & (fsm_output[9]);
  assign and_981_nl = and_dcpl_186 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_983_nl = and_dcpl_171 & and_dcpl_97 & (fsm_output[9]);
  assign and_985_nl = or_dcpl_332 & (fsm_output[9]);
  assign and_990_nl = and_dcpl_183 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_992_nl = and_dcpl_175 & and_dcpl_159 & (fsm_output[9]);
  assign and_994_nl = or_dcpl_334 & (fsm_output[9]);
  assign and_999_nl = and_dcpl_180 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_1001_nl = and_dcpl_175 & and_dcpl_84 & (fsm_output[9]);
  assign and_1003_nl = or_dcpl_336 & (fsm_output[9]);
  assign and_1008_nl = and_dcpl_177 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_1010_nl = and_dcpl_171 & and_dcpl_154 & (fsm_output[9]);
  assign and_1012_nl = or_dcpl_338 & (fsm_output[9]);
  assign and_1017_nl = and_dcpl_173 & (~ LOOPK1_slc_cnt_5_0_66_itm) & (fsm_output[4]);
  assign and_1019_nl = and_dcpl_175 & and_dcpl_97 & (fsm_output[9]);
  assign and_1021_nl = or_dcpl_340 & (fsm_output[9]);
  assign and_1026_nl = and_dcpl_169 & LOOPK1_slc_cnt_5_0_66_itm & (fsm_output[4]);
  assign and_1028_nl = and_dcpl_171 & and_dcpl_159 & (fsm_output[9]);
  assign and_1030_nl = or_dcpl_342 & (fsm_output[9]);
  assign and_1035_nl = and_dcpl_116 & and_dcpl_211 & (fsm_output[4]);
  assign and_1037_nl = and_dcpl_143 & and_dcpl_101 & (fsm_output[9]);
  assign and_1039_nl = or_dcpl_345 & (fsm_output[9]);
  assign and_1044_nl = and_dcpl_122 & and_dcpl_214 & (fsm_output[4]);
  assign and_1046_nl = and_dcpl_139 & and_dcpl_125 & (fsm_output[9]);
  assign and_1048_nl = or_dcpl_348 & (fsm_output[9]);
  assign and_1053_nl = and_dcpl_129 & and_dcpl_211 & (fsm_output[4]);
  assign and_1055_nl = and_dcpl_143 & and_dcpl_91 & (fsm_output[9]);
  assign and_1057_nl = or_dcpl_350 & (fsm_output[9]);
  assign and_1062_nl = and_dcpl_132 & and_dcpl_214 & (fsm_output[4]);
  assign and_1064_nl = and_dcpl_139 & and_dcpl_135 & (fsm_output[9]);
  assign and_1066_nl = or_dcpl_352 & (fsm_output[9]);
  assign and_1071_nl = and_dcpl_137 & and_dcpl_211 & (fsm_output[4]);
  assign and_1073_nl = and_dcpl_127 & and_dcpl_101 & (fsm_output[9]);
  assign and_1075_nl = or_dcpl_354 & (fsm_output[9]);
  assign and_1080_nl = and_dcpl_141 & and_dcpl_214 & (fsm_output[4]);
  assign and_1082_nl = and_dcpl_119 & and_dcpl_125 & (fsm_output[9]);
  assign and_1084_nl = or_dcpl_356 & (fsm_output[9]);
  assign and_1089_nl = and_dcpl_145 & and_dcpl_211 & (fsm_output[4]);
  assign and_1091_nl = and_dcpl_127 & and_dcpl_91 & (fsm_output[9]);
  assign and_1093_nl = or_dcpl_358 & (fsm_output[9]);
  assign and_1098_nl = and_dcpl_148 & and_dcpl_214 & (fsm_output[4]);
  assign and_1100_nl = and_dcpl_119 & and_dcpl_135 & (fsm_output[9]);
  assign and_1102_nl = or_dcpl_360 & (fsm_output[9]);
  assign and_1107_nl = and_dcpl_148 & and_dcpl_211 & (fsm_output[4]);
  assign and_1109_nl = and_dcpl_143 & and_dcpl_84 & (fsm_output[9]);
  assign and_1111_nl = or_dcpl_362 & (fsm_output[9]);
  assign and_1116_nl = and_dcpl_145 & and_dcpl_214 & (fsm_output[4]);
  assign and_1118_nl = and_dcpl_139 & and_dcpl_154 & (fsm_output[9]);
  assign and_1120_nl = or_dcpl_364 & (fsm_output[9]);
  assign and_1125_nl = and_dcpl_141 & and_dcpl_211 & (fsm_output[4]);
  assign and_1127_nl = and_dcpl_143 & and_dcpl_97 & (fsm_output[9]);
  assign and_1129_nl = or_dcpl_366 & (fsm_output[9]);
  assign and_1134_nl = and_dcpl_137 & and_dcpl_214 & (fsm_output[4]);
  assign and_1136_nl = and_dcpl_139 & and_dcpl_159 & (fsm_output[9]);
  assign and_1138_nl = or_dcpl_368 & (fsm_output[9]);
  assign and_1143_nl = and_dcpl_132 & and_dcpl_211 & (fsm_output[4]);
  assign and_1145_nl = and_dcpl_127 & and_dcpl_84 & (fsm_output[9]);
  assign and_1147_nl = or_dcpl_370 & (fsm_output[9]);
  assign and_1152_nl = and_dcpl_129 & and_dcpl_214 & (fsm_output[4]);
  assign and_1154_nl = and_dcpl_119 & and_dcpl_154 & (fsm_output[9]);
  assign and_1156_nl = or_dcpl_372 & (fsm_output[9]);
  assign and_1161_nl = and_dcpl_122 & and_dcpl_211 & (fsm_output[4]);
  assign and_1163_nl = and_dcpl_127 & and_dcpl_97 & (fsm_output[9]);
  assign and_1165_nl = or_dcpl_374 & (fsm_output[9]);
  assign and_1170_nl = and_dcpl_116 & and_dcpl_214 & (fsm_output[4]);
  assign and_1172_nl = and_dcpl_119 & and_dcpl_159 & (fsm_output[9]);
  assign and_1174_nl = or_dcpl_376 & (fsm_output[9]);
  assign LOOPK3_and_60_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_32_lpi_3,
      LOOPK3_exs_126_0);
  assign and_1178_nl = and_dcpl_248 & and_dcpl_246 & (fsm_output[10]);
  assign nor_144_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_759));
  assign or_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0000);
  assign mux_nl = MUX_s_1_2_2(nor_144_nl, or_tmp_759, or_nl);
  assign LOOPK3_and_61_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_30_lpi_3,
      LOOPK3_exs_124_0);
  assign and_1185_nl = and_dcpl_254 & and_dcpl_252 & (fsm_output[10]);
  assign LOOPK3_and_62_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_34_lpi_3,
      LOOPK3_exs_122_0);
  assign and_1192_nl = and_dcpl_256 & and_dcpl_246 & (fsm_output[10]);
  assign nor_145_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_766));
  assign or_1275_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0001);
  assign mux_6_nl = MUX_s_1_2_2(nor_145_nl, or_tmp_766, or_1275_nl);
  assign LOOPK3_and_63_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_28_lpi_3,
      LOOPK3_exs_120_0);
  assign and_1199_nl = and_dcpl_258 & and_dcpl_252 & (fsm_output[10]);
  assign LOOPK3_and_64_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_36_lpi_3,
      LOOPK3_exs_118_0);
  assign and_1206_nl = and_dcpl_258 & and_dcpl_246 & (fsm_output[10]);
  assign nor_146_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_773));
  assign or_1282_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0010);
  assign mux_7_nl = MUX_s_1_2_2(nor_146_nl, or_tmp_773, or_1282_nl);
  assign LOOPK3_and_65_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_26_lpi_3,
      LOOPK3_exs_116_0);
  assign and_1213_nl = and_dcpl_256 & and_dcpl_252 & (fsm_output[10]);
  assign LOOPK3_and_66_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_38_lpi_3,
      LOOPK3_exs_114_0);
  assign and_1220_nl = and_dcpl_254 & and_dcpl_246 & (fsm_output[10]);
  assign nor_147_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_780));
  assign or_1289_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0011);
  assign mux_8_nl = MUX_s_1_2_2(nor_147_nl, or_tmp_780, or_1289_nl);
  assign LOOPK3_and_67_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_24_lpi_3,
      LOOPK3_exs_112_0);
  assign and_1227_nl = and_dcpl_248 & and_dcpl_252 & (fsm_output[10]);
  assign LOOPK3_and_68_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_40_lpi_3,
      LOOPK3_exs_110_0);
  assign and_1234_nl = and_dcpl_248 & and_dcpl_265 & (fsm_output[10]);
  assign nor_148_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_787));
  assign or_1296_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0100);
  assign mux_9_nl = MUX_s_1_2_2(nor_148_nl, or_tmp_787, or_1296_nl);
  assign LOOPK3_and_69_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_22_lpi_3,
      LOOPK3_exs_108_0);
  assign and_1241_nl = and_dcpl_254 & and_dcpl_268 & (fsm_output[10]);
  assign LOOPK3_and_70_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_42_lpi_3,
      LOOPK3_exs_106_0);
  assign and_1248_nl = and_dcpl_256 & and_dcpl_265 & (fsm_output[10]);
  assign nor_149_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_794));
  assign or_1303_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0101);
  assign mux_10_nl = MUX_s_1_2_2(nor_149_nl, or_tmp_794, or_1303_nl);
  assign LOOPK3_and_71_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_20_lpi_3,
      LOOPK3_exs_104_0);
  assign and_1255_nl = and_dcpl_258 & and_dcpl_268 & (fsm_output[10]);
  assign LOOPK3_and_72_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_44_lpi_3,
      LOOPK3_exs_102_0);
  assign and_1262_nl = and_dcpl_258 & and_dcpl_265 & (fsm_output[10]);
  assign nor_150_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_801));
  assign or_1310_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[3:0]!=4'b0110);
  assign mux_11_nl = MUX_s_1_2_2(nor_150_nl, or_tmp_801, or_1310_nl);
  assign LOOPK3_and_73_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_18_lpi_3,
      LOOPK3_exs_100_0);
  assign and_1269_nl = and_dcpl_256 & and_dcpl_268 & (fsm_output[10]);
  assign LOOPK3_and_74_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_46_lpi_3,
      LOOPK3_exs_98_0);
  assign and_1276_nl = and_dcpl_254 & and_dcpl_265 & (fsm_output[10]);
  assign nor_151_nl = ~((LOOPK5_k_sva_5_0[4]) | (~ or_tmp_808));
  assign mux_12_nl = MUX_s_1_2_2(nor_151_nl, or_tmp_808, nand_31_cse);
  assign LOOPK3_and_75_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_16_lpi_3,
      LOOPK3_exs_96_0);
  assign and_1283_nl = and_dcpl_248 & and_dcpl_268 & (fsm_output[10]);
  assign LOOPK3_and_76_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_48_lpi_3,
      LOOPK3_exs_94_0);
  assign and_1290_nl = and_dcpl_248 & and_dcpl_276 & (fsm_output[10]);
  assign and_2736_nl = nand_34_cse & or_tmp_815;
  assign or_1324_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b000);
  assign mux_13_nl = MUX_s_1_2_2(and_2736_nl, or_tmp_815, or_1324_nl);
  assign LOOPK3_and_77_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_14_lpi_3,
      LOOPK3_exs_92_0);
  assign and_1297_nl = and_dcpl_254 & and_dcpl_278 & (fsm_output[10]);
  assign LOOPK3_and_78_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_50_lpi_3,
      LOOPK3_exs_90_0);
  assign and_1304_nl = and_dcpl_256 & and_dcpl_276 & (fsm_output[10]);
  assign and_2738_nl = nand_34_cse & or_tmp_822;
  assign or_1331_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b001);
  assign mux_14_nl = MUX_s_1_2_2(and_2738_nl, or_tmp_822, or_1331_nl);
  assign LOOPK3_and_79_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_12_lpi_3,
      LOOPK3_exs_88_0);
  assign and_1311_nl = and_dcpl_258 & and_dcpl_278 & (fsm_output[10]);
  assign LOOPK3_and_80_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_52_lpi_3,
      LOOPK3_exs_86_0);
  assign and_1318_nl = and_dcpl_258 & and_dcpl_276 & (fsm_output[10]);
  assign and_2740_nl = nand_34_cse & or_tmp_829;
  assign or_1338_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[2:0]!=3'b010);
  assign mux_15_nl = MUX_s_1_2_2(and_2740_nl, or_tmp_829, or_1338_nl);
  assign LOOPK3_and_81_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_10_lpi_3,
      LOOPK3_exs_84_0);
  assign and_1325_nl = and_dcpl_256 & and_dcpl_278 & (fsm_output[10]);
  assign LOOPK3_and_82_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_54_lpi_3,
      LOOPK3_exs_82_0);
  assign and_1332_nl = and_dcpl_254 & and_dcpl_276 & (fsm_output[10]);
  assign and_2742_nl = nand_34_cse & or_tmp_836;
  assign mux_16_nl = MUX_s_1_2_2(and_2742_nl, or_tmp_836, nand_44_cse);
  assign LOOPK3_and_83_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_8_lpi_3,
      LOOPK3_exs_80_0);
  assign and_1339_nl = and_dcpl_248 & and_dcpl_278 & (fsm_output[10]);
  assign LOOPK3_and_84_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_56_lpi_3,
      LOOPK3_exs_78_0);
  assign and_1346_nl = and_dcpl_248 & and_dcpl_286 & (fsm_output[10]);
  assign and_2744_nl = nand_47_cse & or_tmp_843;
  assign or_1352_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[1:0]!=2'b00);
  assign mux_17_nl = MUX_s_1_2_2(and_2744_nl, or_tmp_843, or_1352_nl);
  assign LOOPK3_and_85_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_6_lpi_3,
      LOOPK3_exs_76_0);
  assign and_1353_nl = and_dcpl_254 & and_dcpl_288 & (fsm_output[10]);
  assign LOOPK3_and_86_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_58_lpi_3,
      LOOPK3_exs_74_0);
  assign and_1360_nl = and_dcpl_256 & and_dcpl_286 & (fsm_output[10]);
  assign and_2746_nl = nand_47_cse & or_tmp_850;
  assign or_1359_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[1:0]!=2'b01);
  assign mux_18_nl = MUX_s_1_2_2(and_2746_nl, or_tmp_850, or_1359_nl);
  assign LOOPK3_and_87_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_4_lpi_3,
      LOOPK3_exs_72_0);
  assign and_1367_nl = and_dcpl_258 & and_dcpl_288 & (fsm_output[10]);
  assign LOOPK3_and_88_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_60_lpi_3,
      LOOPK3_exs_70_0);
  assign and_1374_nl = and_dcpl_258 & and_dcpl_286 & (fsm_output[10]);
  assign and_2748_nl = (~((LOOPK5_k_sva_5_0[4:1]==4'b1111))) & or_tmp_857;
  assign or_1366_nl = (~ (fsm_output[7])) | (LOOPK5_k_sva_5_0[0]);
  assign mux_19_nl = MUX_s_1_2_2(and_2748_nl, or_tmp_857, or_1366_nl);
  assign LOOPK3_and_89_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_2_lpi_3,
      LOOPK3_exs_68_0);
  assign and_1381_nl = and_dcpl_256 & and_dcpl_288 & (fsm_output[10]);
  assign LOOPK3_and_90_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_62_lpi_3,
      LOOPK3_exs_66_0);
  assign and_1388_nl = and_dcpl_254 & and_dcpl_286 & (fsm_output[10]);
  assign LOOPK3_and_152_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_31_lpi_3,
      LOOPK3_exs_124_0);
  assign and_1395_nl = and_dcpl_296 & and_dcpl_252 & (fsm_output[10]);
  assign nor_153_nl = ~((fsm_output[10]) | (~ or_tmp_868));
  assign nand_56_nl = ~((LOOPL2_l_sva[5:0]==6'b011111));
  assign mux_20_nl = MUX_s_1_2_2(nor_153_nl, or_tmp_868, nand_56_nl);
  assign LOOPK3_and_153_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_33_lpi_3,
      LOOPK3_exs_126_0);
  assign and_1402_nl = and_dcpl_301 & and_dcpl_246 & (fsm_output[10]);
  assign and_2752_nl = nand_58_cse & or_tmp_873;
  assign or_1381_nl = (LOOPL2_l_sva[4:0]!=5'b00001);
  assign mux_21_nl = MUX_s_1_2_2(and_2752_nl, or_tmp_873, or_1381_nl);
  assign LOOPK3_and_154_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_29_lpi_3,
      LOOPK3_exs_120_0);
  assign and_1409_nl = and_dcpl_303 & and_dcpl_252 & (fsm_output[10]);
  assign nor_154_nl = ~((fsm_output[10]) | (~ or_tmp_878));
  assign or_1386_nl = (LOOPL2_l_sva[5:0]!=6'b011101);
  assign mux_22_nl = MUX_s_1_2_2(nor_154_nl, or_tmp_878, or_1386_nl);
  assign LOOPK3_and_155_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_35_lpi_3,
      LOOPK3_exs_122_0);
  assign and_1416_nl = and_dcpl_305 & and_dcpl_246 & (fsm_output[10]);
  assign and_2754_nl = nand_58_cse & or_tmp_883;
  assign or_1391_nl = (LOOPL2_l_sva[4:0]!=5'b00011);
  assign mux_23_nl = MUX_s_1_2_2(and_2754_nl, or_tmp_883, or_1391_nl);
  assign LOOPK3_and_156_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_27_lpi_3,
      LOOPK3_exs_116_0);
  assign and_1423_nl = and_dcpl_305 & and_dcpl_252 & (fsm_output[10]);
  assign nor_155_nl = ~((fsm_output[10]) | (~ or_tmp_888));
  assign or_1396_nl = (LOOPL2_l_sva[5:0]!=6'b011011);
  assign mux_24_nl = MUX_s_1_2_2(nor_155_nl, or_tmp_888, or_1396_nl);
  assign LOOPK3_and_157_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_37_lpi_3,
      LOOPK3_exs_118_0);
  assign and_1430_nl = and_dcpl_303 & and_dcpl_246 & (fsm_output[10]);
  assign and_2756_nl = nand_58_cse & or_tmp_893;
  assign or_1401_nl = (LOOPL2_l_sva[4:0]!=5'b00101);
  assign mux_25_nl = MUX_s_1_2_2(and_2756_nl, or_tmp_893, or_1401_nl);
  assign LOOPK3_and_158_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_25_lpi_3,
      LOOPK3_exs_112_0);
  assign and_1437_nl = and_dcpl_301 & and_dcpl_252 & (fsm_output[10]);
  assign nor_156_nl = ~((fsm_output[10]) | (~ or_tmp_898));
  assign or_1406_nl = (LOOPL2_l_sva[5:0]!=6'b011001);
  assign mux_26_nl = MUX_s_1_2_2(nor_156_nl, or_tmp_898, or_1406_nl);
  assign LOOPK3_and_159_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_39_lpi_3,
      LOOPK3_exs_114_0);
  assign and_1444_nl = and_dcpl_296 & and_dcpl_246 & (fsm_output[10]);
  assign and_2758_nl = nand_58_cse & or_tmp_903;
  assign or_1411_nl = (LOOPL2_l_sva[4:0]!=5'b00111);
  assign mux_27_nl = MUX_s_1_2_2(and_2758_nl, or_tmp_903, or_1411_nl);
  assign LOOPK3_and_160_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_23_lpi_3,
      LOOPK3_exs_108_0);
  assign and_1451_nl = and_dcpl_296 & and_dcpl_268 & (fsm_output[10]);
  assign nor_157_nl = ~((fsm_output[10]) | (~ or_tmp_908));
  assign or_1416_nl = (LOOPL2_l_sva[5:0]!=6'b010111);
  assign mux_28_nl = MUX_s_1_2_2(nor_157_nl, or_tmp_908, or_1416_nl);
  assign LOOPK3_and_161_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_41_lpi_3,
      LOOPK3_exs_110_0);
  assign and_1458_nl = and_dcpl_301 & and_dcpl_265 & (fsm_output[10]);
  assign and_2760_nl = nand_58_cse & or_tmp_913;
  assign or_1421_nl = (LOOPL2_l_sva[4:0]!=5'b01001);
  assign mux_29_nl = MUX_s_1_2_2(and_2760_nl, or_tmp_913, or_1421_nl);
  assign LOOPK3_and_162_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_21_lpi_3,
      LOOPK3_exs_104_0);
  assign and_1465_nl = and_dcpl_303 & and_dcpl_268 & (fsm_output[10]);
  assign nor_158_nl = ~((fsm_output[10]) | (~ or_tmp_918));
  assign or_1426_nl = (LOOPL2_l_sva[5:0]!=6'b010101);
  assign mux_30_nl = MUX_s_1_2_2(nor_158_nl, or_tmp_918, or_1426_nl);
  assign LOOPK3_and_163_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_43_lpi_3,
      LOOPK3_exs_106_0);
  assign and_1472_nl = and_dcpl_305 & and_dcpl_265 & (fsm_output[10]);
  assign and_2762_nl = nand_58_cse & or_tmp_923;
  assign or_1431_nl = (LOOPL2_l_sva[4:0]!=5'b01011);
  assign mux_31_nl = MUX_s_1_2_2(and_2762_nl, or_tmp_923, or_1431_nl);
  assign LOOPK3_and_164_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_19_lpi_3,
      LOOPK3_exs_100_0);
  assign and_1479_nl = and_dcpl_305 & and_dcpl_268 & (fsm_output[10]);
  assign nor_159_nl = ~((fsm_output[10]) | (~ or_tmp_928));
  assign or_1436_nl = (LOOPL2_l_sva[5:0]!=6'b010011);
  assign mux_32_nl = MUX_s_1_2_2(nor_159_nl, or_tmp_928, or_1436_nl);
  assign LOOPK3_and_165_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_45_lpi_3,
      LOOPK3_exs_102_0);
  assign and_1486_nl = and_dcpl_303 & and_dcpl_265 & (fsm_output[10]);
  assign and_2764_nl = nand_58_cse & or_tmp_933;
  assign or_1441_nl = (LOOPL2_l_sva[4:0]!=5'b01101);
  assign mux_33_nl = MUX_s_1_2_2(and_2764_nl, or_tmp_933, or_1441_nl);
  assign LOOPK3_and_166_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_17_lpi_3,
      LOOPK3_exs_96_0);
  assign and_1493_nl = and_dcpl_301 & and_dcpl_268 & (fsm_output[10]);
  assign nor_160_nl = ~((fsm_output[10]) | (~ or_tmp_938));
  assign or_1446_nl = (LOOPL2_l_sva[5:0]!=6'b010001);
  assign mux_34_nl = MUX_s_1_2_2(nor_160_nl, or_tmp_938, or_1446_nl);
  assign LOOPK3_and_167_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_47_lpi_3,
      LOOPK3_exs_98_0);
  assign and_1500_nl = and_dcpl_296 & and_dcpl_265 & (fsm_output[10]);
  assign and_2766_nl = nand_58_cse & or_tmp_943;
  assign nand_73_nl = ~((LOOPL2_l_sva[4:0]==5'b01111));
  assign mux_35_nl = MUX_s_1_2_2(and_2766_nl, or_tmp_943, nand_73_nl);
  assign LOOPK3_and_168_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_15_lpi_3,
      LOOPK3_exs_92_0);
  assign and_1507_nl = and_dcpl_296 & and_dcpl_278 & (fsm_output[10]);
  assign nor_161_nl = ~((fsm_output[10]) | (~ or_tmp_948));
  assign or_1456_nl = (LOOPL2_l_sva[5:0]!=6'b001111);
  assign mux_36_nl = MUX_s_1_2_2(nor_161_nl, or_tmp_948, or_1456_nl);
  assign LOOPK3_and_169_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_49_lpi_3,
      LOOPK3_exs_94_0);
  assign and_1514_nl = and_dcpl_301 & and_dcpl_276 & (fsm_output[10]);
  assign and_2768_nl = nand_75_cse & or_tmp_953;
  assign or_1461_nl = (LOOPL2_l_sva[3:0]!=4'b0001);
  assign mux_37_nl = MUX_s_1_2_2(and_2768_nl, or_tmp_953, or_1461_nl);
  assign LOOPK3_and_170_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_13_lpi_3,
      LOOPK3_exs_88_0);
  assign and_1521_nl = and_dcpl_303 & and_dcpl_278 & (fsm_output[10]);
  assign nor_162_nl = ~((fsm_output[10]) | (~ or_tmp_958));
  assign or_1466_nl = (LOOPL2_l_sva[5:0]!=6'b001101);
  assign mux_38_nl = MUX_s_1_2_2(nor_162_nl, or_tmp_958, or_1466_nl);
  assign LOOPK3_and_171_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_51_lpi_3,
      LOOPK3_exs_90_0);
  assign and_1528_nl = and_dcpl_305 & and_dcpl_276 & (fsm_output[10]);
  assign and_2770_nl = nand_75_cse & or_tmp_963;
  assign or_1471_nl = (LOOPL2_l_sva[3:0]!=4'b0011);
  assign mux_39_nl = MUX_s_1_2_2(and_2770_nl, or_tmp_963, or_1471_nl);
  assign LOOPK3_and_172_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_11_lpi_3,
      LOOPK3_exs_84_0);
  assign and_1535_nl = and_dcpl_305 & and_dcpl_278 & (fsm_output[10]);
  assign nor_163_nl = ~((fsm_output[10]) | (~ or_tmp_968));
  assign or_1476_nl = (LOOPL2_l_sva[5:0]!=6'b001011);
  assign mux_40_nl = MUX_s_1_2_2(nor_163_nl, or_tmp_968, or_1476_nl);
  assign LOOPK3_and_173_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_53_lpi_3,
      LOOPK3_exs_86_0);
  assign and_1542_nl = and_dcpl_303 & and_dcpl_276 & (fsm_output[10]);
  assign and_2772_nl = nand_75_cse & or_tmp_973;
  assign or_1481_nl = (LOOPL2_l_sva[3:0]!=4'b0101);
  assign mux_41_nl = MUX_s_1_2_2(and_2772_nl, or_tmp_973, or_1481_nl);
  assign LOOPK3_and_174_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_9_lpi_3,
      LOOPK3_exs_80_0);
  assign and_1549_nl = and_dcpl_301 & and_dcpl_278 & (fsm_output[10]);
  assign nor_164_nl = ~((fsm_output[10]) | (~ or_tmp_978));
  assign or_1486_nl = (LOOPL2_l_sva[5:0]!=6'b001001);
  assign mux_42_nl = MUX_s_1_2_2(nor_164_nl, or_tmp_978, or_1486_nl);
  assign LOOPK3_and_175_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_55_lpi_3,
      LOOPK3_exs_82_0);
  assign and_1556_nl = and_dcpl_296 & and_dcpl_276 & (fsm_output[10]);
  assign and_2774_nl = nand_75_cse & or_tmp_983;
  assign nand_82_nl = ~((LOOPL2_l_sva[3:0]==4'b0111));
  assign mux_43_nl = MUX_s_1_2_2(and_2774_nl, or_tmp_983, nand_82_nl);
  assign LOOPK3_and_176_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_7_lpi_3,
      LOOPK3_exs_76_0);
  assign and_1563_nl = and_dcpl_296 & and_dcpl_288 & (fsm_output[10]);
  assign nor_165_nl = ~((fsm_output[10]) | (~ or_tmp_988));
  assign or_1496_nl = (LOOPL2_l_sva[5:0]!=6'b000111);
  assign mux_44_nl = MUX_s_1_2_2(nor_165_nl, or_tmp_988, or_1496_nl);
  assign LOOPK3_and_177_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_57_lpi_3,
      LOOPK3_exs_78_0);
  assign and_1570_nl = and_dcpl_301 & and_dcpl_286 & (fsm_output[10]);
  assign and_2776_nl = nand_84_cse & or_tmp_993;
  assign or_1501_nl = (LOOPL2_l_sva[2:0]!=3'b001);
  assign mux_45_nl = MUX_s_1_2_2(and_2776_nl, or_tmp_993, or_1501_nl);
  assign LOOPK3_and_178_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_5_lpi_3,
      LOOPK3_exs_72_0);
  assign and_1577_nl = and_dcpl_303 & and_dcpl_288 & (fsm_output[10]);
  assign nor_166_nl = ~((fsm_output[10]) | (~ or_tmp_998));
  assign or_1506_nl = (LOOPL2_l_sva[5:0]!=6'b000101);
  assign mux_46_nl = MUX_s_1_2_2(nor_166_nl, or_tmp_998, or_1506_nl);
  assign LOOPK3_and_179_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_59_lpi_3,
      LOOPK3_exs_74_0);
  assign and_1584_nl = and_dcpl_305 & and_dcpl_286 & (fsm_output[10]);
  assign and_2778_nl = nand_84_cse & or_tmp_1003;
  assign or_1511_nl = (LOOPL2_l_sva[2:0]!=3'b011);
  assign mux_47_nl = MUX_s_1_2_2(and_2778_nl, or_tmp_1003, or_1511_nl);
  assign LOOPK3_and_180_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_3_lpi_3,
      LOOPK3_exs_68_0);
  assign and_1591_nl = and_dcpl_305 & and_dcpl_288 & (fsm_output[10]);
  assign nor_167_nl = ~((fsm_output[10]) | (~ or_tmp_1008));
  assign or_1516_nl = (LOOPL2_l_sva[5:0]!=6'b000011);
  assign mux_48_nl = MUX_s_1_2_2(nor_167_nl, or_tmp_1008, or_1516_nl);
  assign LOOPK3_and_181_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_61_lpi_3,
      LOOPK3_exs_70_0);
  assign and_1598_nl = and_dcpl_303 & and_dcpl_286 & (fsm_output[10]);
  assign and_2780_nl = (~((LOOPL2_l_sva[0]) & (LOOPL2_l_sva[2]) & (LOOPL2_l_sva[3])
      & (LOOPL2_l_sva[4]) & (LOOPL2_l_sva[5]) & (fsm_output[10]))) & or_tmp_1012;
  assign mux_49_nl = MUX_s_1_2_2(and_2780_nl, or_tmp_1012, LOOPL2_l_sva[1]);
  assign data_out_or_63_nl = (fsm_output[8:7]!=2'b00);
  assign nor_402_nl = ~(MUX_v_16_2_2(z_out_3, 16'b1111111111111111, data_out_or_63_nl));
  assign or_1744_nl = ((~ nor_14_cse) & (fsm_output[7])) | and_2155_cse;
  assign LOOPK3_and_183_nl = MUX_v_16_2_2(16'b0000000000000000, data_out_63_lpi_3,
      LOOPK3_exs_66_0);
  assign and_1614_nl = and_dcpl_296 & and_dcpl_286 & (fsm_output[10]);
  assign LOOPK3_if_LOOPK3_if_and_nl = (~((~ LOOPK3_if_equal_tmp) | (z_out_2[7])))
      & (z_out_2[0]);
  assign LOOPK1_endflag_mux1h_2_nl = MUX1HOT_s_1_3_2(LOOPL1_LOOPL1_and_tmp, LOOPK3_if_LOOPK3_if_and_nl,
      nor_169_cse, {(fsm_output[3]) , (fsm_output[7]) , (fsm_output[12])});
  assign LOOPL1_l_LOOPL1_l_mux_nl = MUX_s_1_2_2((z_out_1[6]), LOOPK5_k_sva_6, fsm_output[13]);
  assign nl_LOOPL2_acc_1_nl = LOOPL2_l_sva + 32'b00000000000000000000000000000001;
  assign LOOPL2_acc_1_nl = nl_LOOPL2_acc_1_nl[31:0];
  assign cnt_nor_nl = ~((fsm_output[16]) | (fsm_output[14]) | (fsm_output[13]) |
      (fsm_output[1]) | LOOPI1_i_or_cse | (fsm_output[12]));
  assign or_1232_nl = (nor_169_cse & (fsm_output[3])) | (fsm_output[10:5]!=6'b000000)
      | and_363_cse;
  assign LOOPL1_l_LOOPL1_l_mux_1_nl = MUX_v_6_2_2((z_out_1[5:0]), z_out, or_1232_nl);
  assign and_2822_nl = LOOPK5_k_nor_seb & (~((and_363_cse | nor_169_cse) & (fsm_output[3])))
      & (~(and_dcpl_348 & ((fsm_output[8]) | (fsm_output[6]) | (fsm_output[10]))));
  assign or_1732_nl = (fsm_output[8:5]!=4'b0000);
  assign mux_51_nl = MUX_s_1_2_2((fsm_output[3]), mux_tmp_46, or_1732_nl);
  assign or_1736_nl = (~((~ LOOPK2_if_1_equal_1_tmp) | (z_out_1[8:6]!=3'b000))) |
      mux_tmp_46;
  assign mux_52_nl = MUX_s_1_2_2(mux_51_nl, or_1736_nl, fsm_output[11]);
  assign nl_LOOPL1_acc_nl = LOOPL1_ac_int_cctor_sva + conv_s2s_32_38(z_out_6[31:0]);
  assign LOOPL1_acc_nl = nl_LOOPL1_acc_nl[37:0];
  assign operator_16_false_div_nl = div_16_u17_u16(17'b10000000000000000, LOOPJ1_sum2_1_sva);
  assign LOOPJ1_sum2_mux_nl = MUX_v_16_2_2(z_out_3, operator_16_false_div_nl, fsm_output[6]);
  assign not_370_nl = ~ (fsm_output[3]);
  assign data_out_nand_nl = ~((~((fsm_output[13]) | (fsm_output[12]) | (fsm_output[9])))
      & and_dcpl_348);
  assign or_1746_nl = (fsm_output[5]) | (fsm_output[7]) | (fsm_output[11]);
  assign operator_6_false_3_mux_1_nl = MUX_v_6_2_2(LOOPJ1_j_sva, LOOPK5_k_sva_5_0,
      or_1746_nl);
  assign nl_z_out = operator_6_false_3_mux_1_nl + 6'b000001;
  assign z_out = nl_z_out[5:0];
  assign operator_8_false_operator_8_false_and_1_nl = (cnt_sva[7]) & (~ or_1253_itm);
  assign operator_8_false_mux_3_nl = MUX_s_1_2_2((cnt_sva[6]), LOOPK5_k_sva_6, or_1253_itm);
  assign operator_8_false_mux_4_nl = MUX_v_6_2_2((cnt_sva[5:0]), LOOPK5_k_sva_5_0,
      or_1253_itm);
  assign operator_8_false_operator_8_false_or_1_nl = (fsm_output[5]) | (fsm_output[11]);
  assign nl_z_out_1 = conv_u2u_8_9({operator_8_false_operator_8_false_and_1_nl ,
      operator_8_false_mux_3_nl , operator_8_false_mux_4_nl}) + conv_s2u_2_9({operator_8_false_operator_8_false_or_1_nl
      , 1'b1});
  assign z_out_1 = nl_z_out_1[8:0];
  assign operator_7_false_1_operator_7_false_1_and_1_nl = (dim[6]) & (~ (fsm_output[14]));
  assign operator_7_false_1_mux_2_nl = MUX_v_6_2_2((dim[5:0]), length, fsm_output[14]);
  assign nl_z_out_2 = conv_u2u_7_8({operator_7_false_1_operator_7_false_1_and_1_nl
      , operator_7_false_1_mux_2_nl}) + 8'b11111111;
  assign z_out_2 = nl_z_out_2[7:0];
  assign LOOPK2_mux_172_nl = MUX_v_16_2_2(LOOPJ1_sum2_1_sva, z_out_4, fsm_output[10]);
  assign LOOPK2_LOOPK2_mux_1_nl = MUX_v_16_56_2((sum_array_0_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_1_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_2_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_3_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_4_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_5_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_6_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_7_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_8_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_9_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_10_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_11_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_12_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_13_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_14_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_15_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_16_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_17_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_18_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_19_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_20_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_21_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_22_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_23_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_24_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_25_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_26_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_27_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_28_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_29_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_30_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_31_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_32_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_33_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_34_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_35_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_36_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_37_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_38_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_39_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_40_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_41_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_42_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_43_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_44_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_45_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_46_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_47_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_48_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_49_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_50_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_51_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_52_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_53_lpi_5_dfm_1_mx0w1[15:0]), (sum_array_54_lpi_5_dfm_1_mx0w1[15:0]),
      (sum_array_55_lpi_5_dfm_1_mx0w1[15:0]), LOOPK5_k_sva_5_0);
  assign LOOPK2_mux_173_nl = MUX_v_16_2_2(LOOPK2_LOOPK2_mux_1_nl, (z_out_6[31:16]),
      fsm_output[10]);
  assign nl_z_out_3 = LOOPK2_mux_172_nl + LOOPK2_mux_173_nl;
  assign z_out_3 = nl_z_out_3[15:0];
  assign LOOPL1_mux_66_nl = MUX_s_1_2_2((LOOPL1_mux_1_itm[15]), (z_out_5[15]), fsm_output[10]);
  assign LOOPL1_LOOPL1_and_2_nl = LOOPL1_mux_66_nl & (~ (fsm_output[9]));
  assign LOOPL1_mux1h_4_nl = MUX1HOT_v_16_3_2(LOOPL1_mux_1_itm, LOOPJ1_sum2_1_sva,
      z_out_5, {(fsm_output[3]) , (fsm_output[9]) , (fsm_output[10])});
  assign LOOPL2_LOOPL2_mux_1_nl = MUX_v_32_56_2((sum_array_0_lpi_3[31:0]), (sum_array_1_lpi_3[31:0]),
      (sum_array_2_lpi_3[31:0]), (sum_array_3_lpi_3[31:0]), (sum_array_4_lpi_3[31:0]),
      (sum_array_5_lpi_3[31:0]), (sum_array_6_lpi_3[31:0]), (sum_array_7_lpi_3[31:0]),
      (sum_array_8_lpi_3[31:0]), (sum_array_9_lpi_3[31:0]), (sum_array_10_lpi_3[31:0]),
      (sum_array_11_lpi_3[31:0]), (sum_array_12_lpi_3[31:0]), (sum_array_13_lpi_3[31:0]),
      (sum_array_14_lpi_3[31:0]), (sum_array_15_lpi_3[31:0]), (sum_array_16_lpi_3[31:0]),
      (sum_array_17_lpi_3[31:0]), (sum_array_18_lpi_3[31:0]), (sum_array_19_lpi_3[31:0]),
      (sum_array_20_lpi_3[31:0]), (sum_array_21_lpi_3[31:0]), (sum_array_22_lpi_3[31:0]),
      (sum_array_23_lpi_3[31:0]), (sum_array_24_lpi_3[31:0]), (sum_array_25_lpi_3[31:0]),
      (sum_array_26_lpi_3[31:0]), (sum_array_27_lpi_3[31:0]), (sum_array_28_lpi_3[31:0]),
      (sum_array_29_lpi_3[31:0]), (sum_array_30_lpi_3[31:0]), (sum_array_31_lpi_3[31:0]),
      (sum_array_32_lpi_3[31:0]), (sum_array_33_lpi_3[31:0]), (sum_array_34_lpi_3[31:0]),
      (sum_array_35_lpi_3[31:0]), (sum_array_36_lpi_3[31:0]), (sum_array_37_lpi_3[31:0]),
      (sum_array_38_lpi_3[31:0]), (sum_array_39_lpi_3[31:0]), (sum_array_40_lpi_3[31:0]),
      (sum_array_41_lpi_3[31:0]), (sum_array_42_lpi_3[31:0]), (sum_array_43_lpi_3[31:0]),
      (sum_array_44_lpi_3[31:0]), (sum_array_45_lpi_3[31:0]), (sum_array_46_lpi_3[31:0]),
      (sum_array_47_lpi_3[31:0]), (sum_array_48_lpi_3[31:0]), (sum_array_49_lpi_3[31:0]),
      (sum_array_50_lpi_3[31:0]), (sum_array_51_lpi_3[31:0]), (sum_array_52_lpi_3[31:0]),
      (sum_array_53_lpi_3[31:0]), (sum_array_54_lpi_3[31:0]), (sum_array_55_lpi_3[31:0]),
      LOOPK5_k_sva_5_0);
  assign LOOPL1_mux1h_5_nl = MUX1HOT_v_38_3_2(({{22{z_out_5[15]}}, z_out_5}), LOOPK2_mux_169,
      (signext_38_32(LOOPL2_LOOPL2_mux_1_nl)), {(fsm_output[3]) , (fsm_output[9])
      , (fsm_output[10])});
  assign nl_z_out_6 = $signed(({LOOPL1_LOOPL1_and_2_nl , LOOPL1_mux1h_4_nl})) * $signed(conv_u2s_38_39(LOOPL1_mux1h_5_nl));
  assign z_out_6 = nl_z_out_6[37:0];
  assign z_out_4 = MUX_v_16_64_2(data_out_0_lpi_6, data_out_1_lpi_3, data_out_2_lpi_3,
      data_out_3_lpi_3, data_out_4_lpi_3, data_out_5_lpi_3, data_out_6_lpi_3, data_out_7_lpi_3,
      data_out_8_lpi_3, data_out_9_lpi_3, data_out_10_lpi_3, data_out_11_lpi_3, data_out_12_lpi_3,
      data_out_13_lpi_3, data_out_14_lpi_3, data_out_15_lpi_3, data_out_16_lpi_3,
      data_out_17_lpi_3, data_out_18_lpi_3, data_out_19_lpi_3, data_out_20_lpi_3,
      data_out_21_lpi_3, data_out_22_lpi_3, data_out_23_lpi_3, data_out_24_lpi_3,
      data_out_25_lpi_3, data_out_26_lpi_3, data_out_27_lpi_3, data_out_28_lpi_3,
      data_out_29_lpi_3, data_out_30_lpi_3, data_out_31_lpi_3, data_out_32_lpi_3,
      data_out_33_lpi_3, data_out_34_lpi_3, data_out_35_lpi_3, data_out_36_lpi_3,
      data_out_37_lpi_3, data_out_38_lpi_3, data_out_39_lpi_3, data_out_40_lpi_3,
      data_out_41_lpi_3, data_out_42_lpi_3, data_out_43_lpi_3, data_out_44_lpi_3,
      data_out_45_lpi_3, data_out_46_lpi_3, data_out_47_lpi_3, data_out_48_lpi_3,
      data_out_49_lpi_3, data_out_50_lpi_3, data_out_51_lpi_3, data_out_52_lpi_3,
      data_out_53_lpi_3, data_out_54_lpi_3, data_out_55_lpi_3, data_out_56_lpi_3,
      data_out_57_lpi_3, data_out_58_lpi_3, data_out_59_lpi_3, data_out_60_lpi_3,
      data_out_61_lpi_3, data_out_62_lpi_3, data_out_63_lpi_3, LOOPK5_mux_cse);
  assign z_out_5 = MUX_v_16_64_2((k_channel_data_sva[15:0]), (k_channel_data_sva[31:16]),
      (k_channel_data_sva[47:32]), (k_channel_data_sva[63:48]), (k_channel_data_sva[79:64]),
      (k_channel_data_sva[95:80]), (k_channel_data_sva[111:96]), (k_channel_data_sva[127:112]),
      (k_channel_data_sva[143:128]), (k_channel_data_sva[159:144]), (k_channel_data_sva[175:160]),
      (k_channel_data_sva[191:176]), (k_channel_data_sva[207:192]), (k_channel_data_sva[223:208]),
      (k_channel_data_sva[239:224]), (k_channel_data_sva[255:240]), (k_channel_data_sva[271:256]),
      (k_channel_data_sva[287:272]), (k_channel_data_sva[303:288]), (k_channel_data_sva[319:304]),
      (k_channel_data_sva[335:320]), (k_channel_data_sva[351:336]), (k_channel_data_sva[367:352]),
      (k_channel_data_sva[383:368]), (k_channel_data_sva[399:384]), (k_channel_data_sva[415:400]),
      (k_channel_data_sva[431:416]), (k_channel_data_sva[447:432]), (k_channel_data_sva[463:448]),
      (k_channel_data_sva[479:464]), (k_channel_data_sva[495:480]), (k_channel_data_sva[511:496]),
      (k_channel_data_sva[527:512]), (k_channel_data_sva[543:528]), (k_channel_data_sva[559:544]),
      (k_channel_data_sva[575:560]), (k_channel_data_sva[591:576]), (k_channel_data_sva[607:592]),
      (k_channel_data_sva[623:608]), (k_channel_data_sva[639:624]), (k_channel_data_sva[655:640]),
      (k_channel_data_sva[671:656]), (k_channel_data_sva[687:672]), (k_channel_data_sva[703:688]),
      (k_channel_data_sva[719:704]), (k_channel_data_sva[735:720]), (k_channel_data_sva[751:736]),
      (k_channel_data_sva[767:752]), (k_channel_data_sva[783:768]), (k_channel_data_sva[799:784]),
      (k_channel_data_sva[815:800]), (k_channel_data_sva[831:816]), (k_channel_data_sva[847:832]),
      (k_channel_data_sva[863:848]), (k_channel_data_sva[879:864]), (k_channel_data_sva[895:880]),
      (k_channel_data_sva[911:896]), (k_channel_data_sva[927:912]), (k_channel_data_sva[943:928]),
      (k_channel_data_sva[959:944]), (k_channel_data_sva[975:960]), (k_channel_data_sva[991:976]),
      (k_channel_data_sva[1007:992]), (k_channel_data_sva[1023:1008]), LOOPK5_mux_cse);

  function automatic [15:0] div_16_u17_u16;
    input [16:0] l;
    input [15:0] r;
    reg [16:0] rdiv;
    reg [16:0] diff;
    reg [17:0] diff_tmp;
    reg [32:0] lbuf;
    integer i; 
  begin
    lbuf = 33'b0;
    lbuf[16:0] = l;
    for(i=16; i>=0; i=i-1)
    begin
      diff_tmp = (lbuf[32:16] - {1'b0,r});
      diff = diff_tmp[16:0];
      rdiv[i] = ~diff[16];
      if(diff[16] == 0)
        lbuf[32:16] = diff;
      lbuf[32:1] = lbuf[31:0];
    end
    div_16_u17_u16 = rdiv[15:0];
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_3_2;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [2:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    MUX1HOT_v_16_3_2 = result;
  end
  endfunction


  function automatic [37:0] MUX1HOT_v_38_20_2;
    input [37:0] input_19;
    input [37:0] input_18;
    input [37:0] input_17;
    input [37:0] input_16;
    input [37:0] input_15;
    input [37:0] input_14;
    input [37:0] input_13;
    input [37:0] input_12;
    input [37:0] input_11;
    input [37:0] input_10;
    input [37:0] input_9;
    input [37:0] input_8;
    input [37:0] input_7;
    input [37:0] input_6;
    input [37:0] input_5;
    input [37:0] input_4;
    input [37:0] input_3;
    input [37:0] input_2;
    input [37:0] input_1;
    input [37:0] input_0;
    input [19:0] sel;
    reg [37:0] result;
  begin
    result = input_0 & {38{sel[0]}};
    result = result | (input_1 & {38{sel[1]}});
    result = result | (input_2 & {38{sel[2]}});
    result = result | (input_3 & {38{sel[3]}});
    result = result | (input_4 & {38{sel[4]}});
    result = result | (input_5 & {38{sel[5]}});
    result = result | (input_6 & {38{sel[6]}});
    result = result | (input_7 & {38{sel[7]}});
    result = result | (input_8 & {38{sel[8]}});
    result = result | (input_9 & {38{sel[9]}});
    result = result | (input_10 & {38{sel[10]}});
    result = result | (input_11 & {38{sel[11]}});
    result = result | (input_12 & {38{sel[12]}});
    result = result | (input_13 & {38{sel[13]}});
    result = result | (input_14 & {38{sel[14]}});
    result = result | (input_15 & {38{sel[15]}});
    result = result | (input_16 & {38{sel[16]}});
    result = result | (input_17 & {38{sel[17]}});
    result = result | (input_18 & {38{sel[18]}});
    result = result | (input_19 & {38{sel[19]}});
    MUX1HOT_v_38_20_2 = result;
  end
  endfunction


  function automatic [37:0] MUX1HOT_v_38_3_2;
    input [37:0] input_2;
    input [37:0] input_1;
    input [37:0] input_0;
    input [2:0] sel;
    reg [37:0] result;
  begin
    result = input_0 & {38{sel[0]}};
    result = result | (input_1 & {38{sel[1]}});
    result = result | (input_2 & {38{sel[2]}});
    MUX1HOT_v_38_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1023:0] MUX_v_1024_2_2;
    input [1023:0] input_0;
    input [1023:0] input_1;
    input  sel;
    reg [1023:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1024_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_56_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [5:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      default : begin
        result = input_55;
      end
    endcase
    MUX_v_16_56_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_64_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [5:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_16_64_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_56_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [31:0] input_3;
    input [31:0] input_4;
    input [31:0] input_5;
    input [31:0] input_6;
    input [31:0] input_7;
    input [31:0] input_8;
    input [31:0] input_9;
    input [31:0] input_10;
    input [31:0] input_11;
    input [31:0] input_12;
    input [31:0] input_13;
    input [31:0] input_14;
    input [31:0] input_15;
    input [31:0] input_16;
    input [31:0] input_17;
    input [31:0] input_18;
    input [31:0] input_19;
    input [31:0] input_20;
    input [31:0] input_21;
    input [31:0] input_22;
    input [31:0] input_23;
    input [31:0] input_24;
    input [31:0] input_25;
    input [31:0] input_26;
    input [31:0] input_27;
    input [31:0] input_28;
    input [31:0] input_29;
    input [31:0] input_30;
    input [31:0] input_31;
    input [31:0] input_32;
    input [31:0] input_33;
    input [31:0] input_34;
    input [31:0] input_35;
    input [31:0] input_36;
    input [31:0] input_37;
    input [31:0] input_38;
    input [31:0] input_39;
    input [31:0] input_40;
    input [31:0] input_41;
    input [31:0] input_42;
    input [31:0] input_43;
    input [31:0] input_44;
    input [31:0] input_45;
    input [31:0] input_46;
    input [31:0] input_47;
    input [31:0] input_48;
    input [31:0] input_49;
    input [31:0] input_50;
    input [31:0] input_51;
    input [31:0] input_52;
    input [31:0] input_53;
    input [31:0] input_54;
    input [31:0] input_55;
    input [5:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      default : begin
        result = input_55;
      end
    endcase
    MUX_v_32_56_2 = result;
  end
  endfunction


  function automatic [35:0] MUX_v_36_56_2;
    input [35:0] input_0;
    input [35:0] input_1;
    input [35:0] input_2;
    input [35:0] input_3;
    input [35:0] input_4;
    input [35:0] input_5;
    input [35:0] input_6;
    input [35:0] input_7;
    input [35:0] input_8;
    input [35:0] input_9;
    input [35:0] input_10;
    input [35:0] input_11;
    input [35:0] input_12;
    input [35:0] input_13;
    input [35:0] input_14;
    input [35:0] input_15;
    input [35:0] input_16;
    input [35:0] input_17;
    input [35:0] input_18;
    input [35:0] input_19;
    input [35:0] input_20;
    input [35:0] input_21;
    input [35:0] input_22;
    input [35:0] input_23;
    input [35:0] input_24;
    input [35:0] input_25;
    input [35:0] input_26;
    input [35:0] input_27;
    input [35:0] input_28;
    input [35:0] input_29;
    input [35:0] input_30;
    input [35:0] input_31;
    input [35:0] input_32;
    input [35:0] input_33;
    input [35:0] input_34;
    input [35:0] input_35;
    input [35:0] input_36;
    input [35:0] input_37;
    input [35:0] input_38;
    input [35:0] input_39;
    input [35:0] input_40;
    input [35:0] input_41;
    input [35:0] input_42;
    input [35:0] input_43;
    input [35:0] input_44;
    input [35:0] input_45;
    input [35:0] input_46;
    input [35:0] input_47;
    input [35:0] input_48;
    input [35:0] input_49;
    input [35:0] input_50;
    input [35:0] input_51;
    input [35:0] input_52;
    input [35:0] input_53;
    input [35:0] input_54;
    input [35:0] input_55;
    input [5:0] sel;
    reg [35:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      default : begin
        result = input_55;
      end
    endcase
    MUX_v_36_56_2 = result;
  end
  endfunction


  function automatic [37:0] MUX_v_38_2_2;
    input [37:0] input_0;
    input [37:0] input_1;
    input  sel;
    reg [37:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_38_2_2 = result;
  end
  endfunction


  function automatic [37:0] MUX_v_38_56_2;
    input [37:0] input_0;
    input [37:0] input_1;
    input [37:0] input_2;
    input [37:0] input_3;
    input [37:0] input_4;
    input [37:0] input_5;
    input [37:0] input_6;
    input [37:0] input_7;
    input [37:0] input_8;
    input [37:0] input_9;
    input [37:0] input_10;
    input [37:0] input_11;
    input [37:0] input_12;
    input [37:0] input_13;
    input [37:0] input_14;
    input [37:0] input_15;
    input [37:0] input_16;
    input [37:0] input_17;
    input [37:0] input_18;
    input [37:0] input_19;
    input [37:0] input_20;
    input [37:0] input_21;
    input [37:0] input_22;
    input [37:0] input_23;
    input [37:0] input_24;
    input [37:0] input_25;
    input [37:0] input_26;
    input [37:0] input_27;
    input [37:0] input_28;
    input [37:0] input_29;
    input [37:0] input_30;
    input [37:0] input_31;
    input [37:0] input_32;
    input [37:0] input_33;
    input [37:0] input_34;
    input [37:0] input_35;
    input [37:0] input_36;
    input [37:0] input_37;
    input [37:0] input_38;
    input [37:0] input_39;
    input [37:0] input_40;
    input [37:0] input_41;
    input [37:0] input_42;
    input [37:0] input_43;
    input [37:0] input_44;
    input [37:0] input_45;
    input [37:0] input_46;
    input [37:0] input_47;
    input [37:0] input_48;
    input [37:0] input_49;
    input [37:0] input_50;
    input [37:0] input_51;
    input [37:0] input_52;
    input [37:0] input_53;
    input [37:0] input_54;
    input [37:0] input_55;
    input [5:0] sel;
    reg [37:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      default : begin
        result = input_55;
      end
    endcase
    MUX_v_38_56_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_37_1_36;
    input [36:0] vector;
    reg [36:0] tmp;
  begin
    tmp = vector >> 36;
    readslicef_37_1_36 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_39_1_38;
    input [38:0] vector;
    reg [38:0] tmp;
  begin
    tmp = vector >> 38;
    readslicef_39_1_38 = tmp[0:0];
  end
  endfunction


  function automatic [37:0] signext_38_13;
    input [12:0] vector;
  begin
    signext_38_13= {{25{vector[12]}}, vector};
  end
  endfunction


  function automatic [37:0] signext_38_32;
    input [31:0] vector;
  begin
    signext_38_32= {{6{vector[31]}}, vector};
  end
  endfunction


  function automatic [31:0] conv_s2s_8_32 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_32 = {{24{vector[7]}}, vector};
  end
  endfunction


  function automatic [37:0] conv_s2s_32_38 ;
    input [31:0]  vector ;
  begin
    conv_s2s_32_38 = {{6{vector[31]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_s2u_2_9 ;
    input [1:0]  vector ;
  begin
    conv_s2u_2_9 = {{7{vector[1]}}, vector};
  end
  endfunction


  function automatic [38:0] conv_s2u_13_39 ;
    input [12:0]  vector ;
  begin
    conv_s2u_13_39 = {{26{vector[12]}}, vector};
  end
  endfunction


  function automatic [36:0] conv_s2u_36_37 ;
    input [35:0]  vector ;
  begin
    conv_s2u_36_37 = {vector[35], vector};
  end
  endfunction


  function automatic [38:0] conv_s2u_38_39 ;
    input [37:0]  vector ;
  begin
    conv_s2u_38_39 = {vector[37], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [38:0] conv_u2s_38_39 ;
    input [37:0]  vector ;
  begin
    conv_u2s_38_39 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2u_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2u_8_9 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Calculator
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Calculator (
  clk, rst, arst_n, head, length, dim, q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy,
      k_chan2_rsc_dat, k_chan2_rsc_vld, k_chan2_rsc_rdy, v_chan2_rsc_dat, v_chan2_rsc_vld,
      v_chan2_rsc_rdy, dout_chan_rsc_dat, dout_chan_rsc_vld, dout_chan_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [1023:0] q_chan2_rsc_dat;
  input q_chan2_rsc_vld;
  output q_chan2_rsc_rdy;
  input [1023:0] k_chan2_rsc_dat;
  input k_chan2_rsc_vld;
  output k_chan2_rsc_rdy;
  input [1023:0] v_chan2_rsc_dat;
  input v_chan2_rsc_vld;
  output v_chan2_rsc_rdy;
  output [15:0] dout_chan_rsc_dat;
  output dout_chan_rsc_vld;
  input dout_chan_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ATTENTION_IP_Attention_Calculator_run ATTENTION_IP_Attention_Calculator_run_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .q_chan2_rsc_dat(q_chan2_rsc_dat),
      .q_chan2_rsc_vld(q_chan2_rsc_vld),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy),
      .k_chan2_rsc_dat(k_chan2_rsc_dat),
      .k_chan2_rsc_vld(k_chan2_rsc_vld),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy),
      .v_chan2_rsc_dat(v_chan2_rsc_dat),
      .v_chan2_rsc_vld(v_chan2_rsc_vld),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy),
      .dout_chan_rsc_dat(dout_chan_rsc_dat),
      .dout_chan_rsc_vld(dout_chan_rsc_vld),
      .dout_chan_rsc_rdy(dout_chan_rsc_rdy)
    );
endmodule




//------> ../ATTENTION_IP_Attention_Filter.v2/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   b08092@cad29.ee.ntu.edu.tw
//  Generated date: Wed Jun 12 20:16:44 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, LOOPI1_C_0_tr0, LOOPK1_C_0_tr0, LOOPL1_C_0_tr0,
      LOOPK2_C_3_tr0, LOOPK3_C_1_tr0, LOOPJ1_C_4_tr0, LOOPI2_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [16:0] fsm_output;
  reg [16:0] fsm_output;
  input LOOPI1_C_0_tr0;
  input LOOPK1_C_0_tr0;
  input LOOPL1_C_0_tr0;
  input LOOPK2_C_3_tr0;
  input LOOPK3_C_1_tr0;
  input LOOPJ1_C_4_tr0;
  input LOOPI2_C_0_tr0;


  // FSM State Type Declaration for ATTENTION_IP_Attention_Filter_run_run_fsm_1
  parameter
    main_C_0 = 5'd0,
    LOOPI1_C_0 = 5'd1,
    LOOPJ1_C_0 = 5'd2,
    LOOPJ1_C_1 = 5'd3,
    LOOPK1_C_0 = 5'd4,
    LOOPJ1_C_2 = 5'd5,
    LOOPK2_C_0 = 5'd6,
    LOOPL1_C_0 = 5'd7,
    LOOPK2_C_1 = 5'd8,
    LOOPK2_C_2 = 5'd9,
    LOOPK2_C_3 = 5'd10,
    LOOPJ1_C_3 = 5'd11,
    LOOPK3_C_0 = 5'd12,
    LOOPK3_C_1 = 5'd13,
    LOOPJ1_C_4 = 5'd14,
    LOOPI2_C_0 = 5'd15,
    main_C_1 = 5'd16;

  reg [4:0] state_var;
  reg [4:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ATTENTION_IP_Attention_Filter_run_run_fsm_1
    case (state_var)
      LOOPI1_C_0 : begin
        fsm_output = 17'b00000000000000010;
        if ( LOOPI1_C_0_tr0 ) begin
          state_var_NS = LOOPJ1_C_0;
        end
        else begin
          state_var_NS = LOOPI1_C_0;
        end
      end
      LOOPJ1_C_0 : begin
        fsm_output = 17'b00000000000000100;
        state_var_NS = LOOPJ1_C_1;
      end
      LOOPJ1_C_1 : begin
        fsm_output = 17'b00000000000001000;
        state_var_NS = LOOPK1_C_0;
      end
      LOOPK1_C_0 : begin
        fsm_output = 17'b00000000000010000;
        if ( LOOPK1_C_0_tr0 ) begin
          state_var_NS = LOOPJ1_C_2;
        end
        else begin
          state_var_NS = LOOPK1_C_0;
        end
      end
      LOOPJ1_C_2 : begin
        fsm_output = 17'b00000000000100000;
        state_var_NS = LOOPK2_C_0;
      end
      LOOPK2_C_0 : begin
        fsm_output = 17'b00000000001000000;
        state_var_NS = LOOPL1_C_0;
      end
      LOOPL1_C_0 : begin
        fsm_output = 17'b00000000010000000;
        if ( LOOPL1_C_0_tr0 ) begin
          state_var_NS = LOOPK2_C_1;
        end
        else begin
          state_var_NS = LOOPL1_C_0;
        end
      end
      LOOPK2_C_1 : begin
        fsm_output = 17'b00000000100000000;
        state_var_NS = LOOPK2_C_2;
      end
      LOOPK2_C_2 : begin
        fsm_output = 17'b00000001000000000;
        state_var_NS = LOOPK2_C_3;
      end
      LOOPK2_C_3 : begin
        fsm_output = 17'b00000010000000000;
        if ( LOOPK2_C_3_tr0 ) begin
          state_var_NS = LOOPJ1_C_3;
        end
        else begin
          state_var_NS = LOOPK2_C_0;
        end
      end
      LOOPJ1_C_3 : begin
        fsm_output = 17'b00000100000000000;
        state_var_NS = LOOPK3_C_0;
      end
      LOOPK3_C_0 : begin
        fsm_output = 17'b00001000000000000;
        state_var_NS = LOOPK3_C_1;
      end
      LOOPK3_C_1 : begin
        fsm_output = 17'b00010000000000000;
        if ( LOOPK3_C_1_tr0 ) begin
          state_var_NS = LOOPJ1_C_4;
        end
        else begin
          state_var_NS = LOOPK3_C_0;
        end
      end
      LOOPJ1_C_4 : begin
        fsm_output = 17'b00100000000000000;
        if ( LOOPJ1_C_4_tr0 ) begin
          state_var_NS = LOOPI2_C_0;
        end
        else begin
          state_var_NS = LOOPJ1_C_0;
        end
      end
      LOOPI2_C_0 : begin
        fsm_output = 17'b01000000000000000;
        if ( LOOPI2_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = LOOPJ1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 17'b10000000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 17'b00000000000000001;
        state_var_NS = LOOPI1_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_staller
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_staller (
  run_wen, q_chan1_rsci_wen_comp, k_chan1_rsci_wen_comp, v_chan1_rsci_wen_comp, q_chan2_rsci_wen_comp,
      k_chan2_rsci_wen_comp, v_chan2_rsci_wen_comp
);
  output run_wen;
  input q_chan1_rsci_wen_comp;
  input k_chan1_rsci_wen_comp;
  input v_chan1_rsci_wen_comp;
  input q_chan2_rsci_wen_comp;
  input k_chan2_rsci_wen_comp;
  input v_chan2_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = q_chan1_rsci_wen_comp & k_chan1_rsci_wen_comp & v_chan1_rsci_wen_comp
      & q_chan2_rsci_wen_comp & k_chan2_rsci_wen_comp & v_chan2_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_v_chan2_rsci_v_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_v_chan2_rsci_v_chan2_wait_ctrl (
  v_chan2_rsci_iswt0, v_chan2_rsci_biwt, v_chan2_rsci_irdy
);
  input v_chan2_rsci_iswt0;
  output v_chan2_rsci_biwt;
  input v_chan2_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign v_chan2_rsci_biwt = v_chan2_rsci_iswt0 & v_chan2_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_k_chan2_rsci_k_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_k_chan2_rsci_k_chan2_wait_ctrl (
  k_chan2_rsci_iswt0, k_chan2_rsci_biwt, k_chan2_rsci_irdy
);
  input k_chan2_rsci_iswt0;
  output k_chan2_rsci_biwt;
  input k_chan2_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign k_chan2_rsci_biwt = k_chan2_rsci_iswt0 & k_chan2_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_q_chan2_rsci_q_chan2_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_q_chan2_rsci_q_chan2_wait_ctrl (
  q_chan2_rsci_iswt0, q_chan2_rsci_biwt, q_chan2_rsci_irdy
);
  input q_chan2_rsci_iswt0;
  output q_chan2_rsci_biwt;
  input q_chan2_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign q_chan2_rsci_biwt = q_chan2_rsci_iswt0 & q_chan2_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_v_chan1_rsci_v_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_v_chan1_rsci_v_chan1_wait_ctrl (
  v_chan1_rsci_iswt0, v_chan1_rsci_biwt, v_chan1_rsci_ivld
);
  input v_chan1_rsci_iswt0;
  output v_chan1_rsci_biwt;
  input v_chan1_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign v_chan1_rsci_biwt = v_chan1_rsci_iswt0 & v_chan1_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_k_chan1_rsci_k_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_k_chan1_rsci_k_chan1_wait_ctrl (
  k_chan1_rsci_iswt0, k_chan1_rsci_biwt, k_chan1_rsci_ivld
);
  input k_chan1_rsci_iswt0;
  output k_chan1_rsci_biwt;
  input k_chan1_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign k_chan1_rsci_biwt = k_chan1_rsci_iswt0 & k_chan1_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_q_chan1_rsci_q_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_q_chan1_rsci_q_chan1_wait_ctrl (
  q_chan1_rsci_iswt0, q_chan1_rsci_biwt, q_chan1_rsci_ivld
);
  input q_chan1_rsci_iswt0;
  output q_chan1_rsci_biwt;
  input q_chan1_rsci_ivld;



  // Interconnect Declarations for Component Instantiations 
  assign q_chan1_rsci_biwt = q_chan1_rsci_iswt0 & q_chan1_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_v_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_v_chan2_rsci (
  v_chan2_rsc_dat, v_chan2_rsc_vld, v_chan2_rsc_rdy, v_chan2_rsci_oswt, v_chan2_rsci_wen_comp,
      v_chan2_rsci_idat
);
  output [1023:0] v_chan2_rsc_dat;
  output v_chan2_rsc_vld;
  input v_chan2_rsc_rdy;
  input v_chan2_rsci_oswt;
  output v_chan2_rsci_wen_comp;
  input [1023:0] v_chan2_rsci_idat;


  // Interconnect Declarations
  wire v_chan2_rsci_biwt;
  wire v_chan2_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd9),
  .width(32'sd1024)) v_chan2_rsci (
      .irdy(v_chan2_rsci_irdy),
      .ivld(v_chan2_rsci_oswt),
      .idat(v_chan2_rsci_idat),
      .rdy(v_chan2_rsc_rdy),
      .vld(v_chan2_rsc_vld),
      .dat(v_chan2_rsc_dat)
    );
  ATTENTION_IP_Attention_Filter_run_v_chan2_rsci_v_chan2_wait_ctrl ATTENTION_IP_Attention_Filter_run_v_chan2_rsci_v_chan2_wait_ctrl_inst
      (
      .v_chan2_rsci_iswt0(v_chan2_rsci_oswt),
      .v_chan2_rsci_biwt(v_chan2_rsci_biwt),
      .v_chan2_rsci_irdy(v_chan2_rsci_irdy)
    );
  assign v_chan2_rsci_wen_comp = (~ v_chan2_rsci_oswt) | v_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_k_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_k_chan2_rsci (
  k_chan2_rsc_dat, k_chan2_rsc_vld, k_chan2_rsc_rdy, k_chan2_rsci_oswt, k_chan2_rsci_wen_comp,
      k_chan2_rsci_idat
);
  output [1023:0] k_chan2_rsc_dat;
  output k_chan2_rsc_vld;
  input k_chan2_rsc_rdy;
  input k_chan2_rsci_oswt;
  output k_chan2_rsci_wen_comp;
  input [1023:0] k_chan2_rsci_idat;


  // Interconnect Declarations
  wire k_chan2_rsci_biwt;
  wire k_chan2_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd8),
  .width(32'sd1024)) k_chan2_rsci (
      .irdy(k_chan2_rsci_irdy),
      .ivld(k_chan2_rsci_oswt),
      .idat(k_chan2_rsci_idat),
      .rdy(k_chan2_rsc_rdy),
      .vld(k_chan2_rsc_vld),
      .dat(k_chan2_rsc_dat)
    );
  ATTENTION_IP_Attention_Filter_run_k_chan2_rsci_k_chan2_wait_ctrl ATTENTION_IP_Attention_Filter_run_k_chan2_rsci_k_chan2_wait_ctrl_inst
      (
      .k_chan2_rsci_iswt0(k_chan2_rsci_oswt),
      .k_chan2_rsci_biwt(k_chan2_rsci_biwt),
      .k_chan2_rsci_irdy(k_chan2_rsci_irdy)
    );
  assign k_chan2_rsci_wen_comp = (~ k_chan2_rsci_oswt) | k_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_q_chan2_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_q_chan2_rsci (
  q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy, q_chan2_rsci_oswt, q_chan2_rsci_wen_comp,
      q_chan2_rsci_idat
);
  output [1023:0] q_chan2_rsc_dat;
  output q_chan2_rsc_vld;
  input q_chan2_rsc_rdy;
  input q_chan2_rsci_oswt;
  output q_chan2_rsci_wen_comp;
  input [1023:0] q_chan2_rsci_idat;


  // Interconnect Declarations
  wire q_chan2_rsci_biwt;
  wire q_chan2_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd7),
  .width(32'sd1024)) q_chan2_rsci (
      .irdy(q_chan2_rsci_irdy),
      .ivld(q_chan2_rsci_oswt),
      .idat(q_chan2_rsci_idat),
      .rdy(q_chan2_rsc_rdy),
      .vld(q_chan2_rsc_vld),
      .dat(q_chan2_rsc_dat)
    );
  ATTENTION_IP_Attention_Filter_run_q_chan2_rsci_q_chan2_wait_ctrl ATTENTION_IP_Attention_Filter_run_q_chan2_rsci_q_chan2_wait_ctrl_inst
      (
      .q_chan2_rsci_iswt0(q_chan2_rsci_oswt),
      .q_chan2_rsci_biwt(q_chan2_rsci_biwt),
      .q_chan2_rsci_irdy(q_chan2_rsci_irdy)
    );
  assign q_chan2_rsci_wen_comp = (~ q_chan2_rsci_oswt) | q_chan2_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_v_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_v_chan1_rsci (
  v_chan1_rsc_dat, v_chan1_rsc_vld, v_chan1_rsc_rdy, v_chan1_rsci_oswt, v_chan1_rsci_wen_comp,
      v_chan1_rsci_idat_mxwt
);
  input [1023:0] v_chan1_rsc_dat;
  input v_chan1_rsc_vld;
  output v_chan1_rsc_rdy;
  input v_chan1_rsci_oswt;
  output v_chan1_rsci_wen_comp;
  output [1023:0] v_chan1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire v_chan1_rsci_biwt;
  wire v_chan1_rsci_ivld;
  wire [1023:0] v_chan1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd6),
  .width(32'sd1024)) v_chan1_rsci (
      .rdy(v_chan1_rsc_rdy),
      .vld(v_chan1_rsc_vld),
      .dat(v_chan1_rsc_dat),
      .irdy(v_chan1_rsci_oswt),
      .ivld(v_chan1_rsci_ivld),
      .idat(v_chan1_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_v_chan1_rsci_v_chan1_wait_ctrl ATTENTION_IP_Attention_Filter_run_v_chan1_rsci_v_chan1_wait_ctrl_inst
      (
      .v_chan1_rsci_iswt0(v_chan1_rsci_oswt),
      .v_chan1_rsci_biwt(v_chan1_rsci_biwt),
      .v_chan1_rsci_ivld(v_chan1_rsci_ivld)
    );
  assign v_chan1_rsci_idat_mxwt = v_chan1_rsci_idat;
  assign v_chan1_rsci_wen_comp = (~ v_chan1_rsci_oswt) | v_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_k_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_k_chan1_rsci (
  k_chan1_rsc_dat, k_chan1_rsc_vld, k_chan1_rsc_rdy, k_chan1_rsci_oswt, k_chan1_rsci_wen_comp,
      k_chan1_rsci_idat_mxwt
);
  input [1023:0] k_chan1_rsc_dat;
  input k_chan1_rsc_vld;
  output k_chan1_rsc_rdy;
  input k_chan1_rsci_oswt;
  output k_chan1_rsci_wen_comp;
  output [1023:0] k_chan1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire k_chan1_rsci_biwt;
  wire k_chan1_rsci_ivld;
  wire [1023:0] k_chan1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd5),
  .width(32'sd1024)) k_chan1_rsci (
      .rdy(k_chan1_rsc_rdy),
      .vld(k_chan1_rsc_vld),
      .dat(k_chan1_rsc_dat),
      .irdy(k_chan1_rsci_oswt),
      .ivld(k_chan1_rsci_ivld),
      .idat(k_chan1_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_k_chan1_rsci_k_chan1_wait_ctrl ATTENTION_IP_Attention_Filter_run_k_chan1_rsci_k_chan1_wait_ctrl_inst
      (
      .k_chan1_rsci_iswt0(k_chan1_rsci_oswt),
      .k_chan1_rsci_biwt(k_chan1_rsci_biwt),
      .k_chan1_rsci_ivld(k_chan1_rsci_ivld)
    );
  assign k_chan1_rsci_idat_mxwt = k_chan1_rsci_idat;
  assign k_chan1_rsci_wen_comp = (~ k_chan1_rsci_oswt) | k_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run_q_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run_q_chan1_rsci (
  q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy, q_chan1_rsci_oswt, q_chan1_rsci_wen_comp,
      q_chan1_rsci_idat_mxwt
);
  input [1023:0] q_chan1_rsc_dat;
  input q_chan1_rsc_vld;
  output q_chan1_rsc_rdy;
  input q_chan1_rsci_oswt;
  output q_chan1_rsci_wen_comp;
  output [1023:0] q_chan1_rsci_idat_mxwt;


  // Interconnect Declarations
  wire q_chan1_rsci_biwt;
  wire q_chan1_rsci_ivld;
  wire [1023:0] q_chan1_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd4),
  .width(32'sd1024)) q_chan1_rsci (
      .rdy(q_chan1_rsc_rdy),
      .vld(q_chan1_rsc_vld),
      .dat(q_chan1_rsc_dat),
      .irdy(q_chan1_rsci_oswt),
      .ivld(q_chan1_rsci_ivld),
      .idat(q_chan1_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_q_chan1_rsci_q_chan1_wait_ctrl ATTENTION_IP_Attention_Filter_run_q_chan1_rsci_q_chan1_wait_ctrl_inst
      (
      .q_chan1_rsci_iswt0(q_chan1_rsci_oswt),
      .q_chan1_rsci_biwt(q_chan1_rsci_biwt),
      .q_chan1_rsci_ivld(q_chan1_rsci_ivld)
    );
  assign q_chan1_rsci_idat_mxwt = q_chan1_rsci_idat;
  assign q_chan1_rsci_wen_comp = (~ q_chan1_rsci_oswt) | q_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter_run
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter_run (
  clk, rst, arst_n, head, length, dim, q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy,
      k_chan1_rsc_dat, k_chan1_rsc_vld, k_chan1_rsc_rdy, v_chan1_rsc_dat, v_chan1_rsc_vld,
      v_chan1_rsc_rdy, q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy, k_chan2_rsc_dat,
      k_chan2_rsc_vld, k_chan2_rsc_rdy, v_chan2_rsc_dat, v_chan2_rsc_vld, v_chan2_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [1023:0] q_chan1_rsc_dat;
  input q_chan1_rsc_vld;
  output q_chan1_rsc_rdy;
  input [1023:0] k_chan1_rsc_dat;
  input k_chan1_rsc_vld;
  output k_chan1_rsc_rdy;
  input [1023:0] v_chan1_rsc_dat;
  input v_chan1_rsc_vld;
  output v_chan1_rsc_rdy;
  output [1023:0] q_chan2_rsc_dat;
  output q_chan2_rsc_vld;
  input q_chan2_rsc_rdy;
  output [1023:0] k_chan2_rsc_dat;
  output k_chan2_rsc_vld;
  input k_chan2_rsc_rdy;
  output [1023:0] v_chan2_rsc_dat;
  output v_chan2_rsc_vld;
  input v_chan2_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire q_chan1_rsci_wen_comp;
  wire [1023:0] q_chan1_rsci_idat_mxwt;
  wire k_chan1_rsci_wen_comp;
  wire [1023:0] k_chan1_rsci_idat_mxwt;
  wire v_chan1_rsci_wen_comp;
  wire [1023:0] v_chan1_rsci_idat_mxwt;
  wire q_chan2_rsci_wen_comp;
  reg [1023:0] q_chan2_rsci_idat;
  wire k_chan2_rsci_wen_comp;
  reg [1023:0] k_chan2_rsci_idat;
  wire v_chan2_rsci_wen_comp;
  reg [1023:0] v_chan2_rsci_idat;
  wire [16:0] fsm_output;
  wire LOOPI2_LOOPI2_if_LOOPI2_if_nor_tmp;
  wire LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp;
  wire LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp;
  wire LOOPK3_if_1_mux_tmp;
  wire LOOPL1_LOOPL1_if_LOOPL1_if_nor_tmp;
  wire LOOPK1_if_unequal_tmp;
  wire LOOPK1_if_equal_tmp;
  wire or_tmp_11;
  wire mux_tmp_3;
  wire or_tmp_198;
  wire and_65_cse;
  wire and_50_cse;
  wire and_52_cse;
  reg LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt;
  reg [19:0] operator_20_true_acc_3_itm_21_2;
  wire [20:0] nl_operator_20_true_acc_3_itm_21_2;
  reg [19:0] avg_sva;
  reg [13:0] max_sva;
  reg reg_q_chan1_rsci_oswt_cse;
  reg reg_k_chan1_rsci_oswt_cse;
  reg reg_v_chan1_rsci_oswt_cse;
  reg reg_q_chan2_rsci_oswt_cse;
  reg reg_k_chan2_rsci_oswt_cse;
  reg reg_v_chan2_rsci_oswt_cse;
  wire sel_and_1_cse;
  wire sel_and_2_cse;
  wire LOOPK2_if_1_LOOPK2_if_1_nor_2_cse;
  reg [5:0] LOOPI1_i_1_6_1_sva;
  wire LOOPL1_l_nand_seb;
  wire and_cse;
  reg [13:0] LOOPK2_mux_106_itm;
  wire LOOPK2_if_1_or_56_itm;
  wire [3:0] z_out;
  wire [4:0] nl_z_out;
  wire [6:0] z_out_1;
  wire [7:0] nl_z_out_1;
  wire [5:0] z_out_2;
  wire [6:0] nl_z_out_2;
  wire [20:0] z_out_3;
  wire [21:0] nl_z_out_3;
  wire [7:0] z_out_4;
  wire [8:0] nl_z_out_4;
  reg [3:0] LOOPI2_i_sva;
  reg sel_28_lpi_3;
  reg sel_26_lpi_3;
  reg sel_30_lpi_3;
  reg sel_24_lpi_3;
  reg sel_32_lpi_3;
  reg sel_22_lpi_3;
  reg sel_34_lpi_3;
  reg sel_20_lpi_3;
  reg sel_36_lpi_3;
  reg sel_18_lpi_3;
  reg sel_38_lpi_3;
  reg sel_16_lpi_3;
  reg sel_40_lpi_3;
  reg sel_14_lpi_3;
  reg sel_42_lpi_3;
  reg sel_12_lpi_3;
  reg sel_44_lpi_3;
  reg sel_10_lpi_3;
  reg sel_46_lpi_3;
  reg sel_8_lpi_3;
  reg sel_48_lpi_3;
  reg sel_6_lpi_3;
  reg sel_50_lpi_3;
  reg sel_4_lpi_3;
  reg sel_52_lpi_3;
  reg sel_2_lpi_3;
  reg sel_54_lpi_3;
  reg sel_27_lpi_3;
  reg sel_29_lpi_3;
  reg sel_25_lpi_3;
  reg sel_31_lpi_3;
  reg sel_23_lpi_3;
  reg sel_33_lpi_3;
  reg sel_21_lpi_3;
  reg sel_35_lpi_3;
  reg sel_19_lpi_3;
  reg sel_37_lpi_3;
  reg sel_17_lpi_3;
  reg sel_39_lpi_3;
  reg sel_15_lpi_3;
  reg sel_41_lpi_3;
  reg sel_13_lpi_3;
  reg sel_43_lpi_3;
  reg sel_11_lpi_3;
  reg sel_45_lpi_3;
  reg sel_9_lpi_3;
  reg sel_47_lpi_3;
  reg sel_7_lpi_3;
  reg sel_49_lpi_3;
  reg sel_5_lpi_3;
  reg sel_51_lpi_3;
  reg sel_3_lpi_3;
  reg sel_53_lpi_3;
  reg sel_1_lpi_3;
  reg sel_55_lpi_3;
  reg [1023:0] q_channel_data_sva;
  reg [1023:0] k_channel_data_sva;
  reg [19:0] LOOPK2_acc_2_itm;
  wire LOOPI1_i_1_6_1_sva_mx0c1;
  wire sel_1_lpi_3_mx0c0;
  wire LOOPK2_k_sva_mx0c1;
  wire LOOPK2_k_sva_mx0c2;
  wire LOOPK1_and_stg_3_1_sva_1;
  wire LOOPK1_and_stg_3_2_sva_1;
  wire LOOPK1_and_stg_3_3_sva_1;
  wire LOOPK1_and_stg_3_4_sva_1;
  wire LOOPK1_and_stg_3_5_sva_1;
  wire LOOPK1_and_stg_3_6_sva_1;
  wire LOOPK1_and_stg_3_7_sva_1;
  wire LOOPK1_and_stg_3_8_sva_1;
  wire LOOPK1_and_stg_3_9_sva_1;
  wire LOOPK1_and_stg_3_10_sva_1;
  wire LOOPK1_and_stg_3_11_sva_1;
  wire LOOPK1_and_stg_2_4_sva_1;
  wire LOOPK1_and_stg_2_5_sva_1;
  wire LOOPK1_and_stg_2_6_sva_1;
  wire LOOPK1_and_stg_2_7_sva_1;
  wire LOOPK1_and_stg_2_0_sva_1;
  wire LOOPK1_and_stg_2_1_sva_1;
  wire LOOPK1_and_stg_2_2_sva_1;
  wire LOOPK1_and_stg_2_3_sva_1;
  wire LOOPK1_and_stg_1_0_sva_1;
  wire LOOPK1_and_stg_1_1_sva_1;
  wire LOOPK1_and_stg_1_2_sva_1;
  wire LOOPK1_and_stg_1_3_sva_1;
  wire LOOPK1_not_127;
  wire LOOPK1_not_129;
  wire LOOPK1_not_131;
  wire LOOPK1_not_133;
  wire LOOPK1_not_135;
  wire LOOPK1_not_137;
  wire LOOPK1_not_139;
  wire LOOPK1_not_141;
  wire LOOPK1_not_143;
  wire LOOPK1_not_145;
  wire LOOPK1_not_147;
  wire LOOPK1_not_149;
  wire LOOPK1_not_151;
  wire LOOPK1_not_153;
  wire LOOPK1_not_155;
  wire LOOPK1_not_157;
  wire LOOPK1_not_159;
  wire LOOPK1_not_161;
  wire LOOPK1_not_163;
  wire LOOPK1_not_165;
  wire LOOPK1_not_167;
  wire LOOPK1_not_169;
  wire LOOPK1_not_171;
  wire LOOPK1_not_173;
  wire LOOPK1_not_175;
  wire LOOPK1_not_177;
  wire LOOPK1_not_179;
  wire LOOPK2_mux_106_itm_mx0c2;
  wire [15:0] operator_16_true_slc_q_channel_data_16_15_0_tmp_sva_1;
  wire [15:0] operator_16_true_1_slc_k_channel_data_16_15_0_tmp_sva_1;
  wire LOOPK2_if_1_and_stg_4_23_sva_1;
  wire LOOPK2_if_1_and_stg_4_22_sva_1;
  wire LOOPK2_if_1_and_stg_4_21_sva_1;
  wire LOOPK2_if_1_and_stg_4_20_sva_1;
  wire LOOPK2_if_1_and_stg_4_19_sva_1;
  wire LOOPK2_if_1_and_stg_4_18_sva_1;
  wire LOOPK2_if_1_and_stg_4_17_sva_1;
  wire LOOPK2_if_1_and_stg_4_16_sva_1;
  wire LOOPK2_if_1_and_stg_4_15_sva_1;
  wire LOOPK2_if_1_and_stg_4_14_sva_1;
  wire LOOPK2_if_1_and_stg_4_13_sva_1;
  wire LOOPK2_if_1_and_stg_4_12_sva_1;
  wire LOOPK2_if_1_and_stg_4_11_sva_1;
  wire LOOPK2_if_1_and_stg_4_10_sva_1;
  wire LOOPK2_if_1_and_stg_4_9_sva_1;
  wire LOOPK2_if_1_and_stg_4_8_sva_1;
  wire LOOPK2_if_1_and_stg_4_7_sva_1;
  wire LOOPK2_if_1_and_stg_4_6_sva_1;
  wire LOOPK2_if_1_and_stg_4_5_sva_1;
  wire LOOPK2_if_1_and_stg_4_4_sva_1;
  wire LOOPK2_if_1_and_stg_4_3_sva_1;
  wire LOOPK2_if_1_and_stg_4_2_sva_1;
  wire LOOPK2_if_1_and_stg_4_1_sva_1;
  wire LOOPK2_if_1_and_stg_3_0_sva_1;
  wire LOOPK2_if_1_and_stg_3_15_sva_1;
  wire LOOPK2_if_1_and_stg_3_14_sva_1;
  wire LOOPK2_if_1_and_stg_3_13_sva_1;
  wire LOOPK2_if_1_and_stg_3_12_sva_1;
  reg LOOPL1_l_sva_6;
  reg [5:0] LOOPL1_l_sva_5_0;
  wire or_7_cse;
  wire LOOPI1_i_LOOPI1_i_LOOPI1_i_nor_cse;
  wire or_282_itm;
  reg LOOPK2_k_sva_rsp_0;
  reg [4:0] LOOPK2_k_sva_rsp_1;
  wire LOOPK2_k_and_ssc;

  wire LOOPK2_if_1_not_nl;
  wire LOOPI1_i_not_nl;
  wire sel_mux_nl;
  wire sel_nand_nl;
  wire sel_nor_nl;
  wire LOOPK1_and_73_nl;
  wire LOOPK2_if_1_or_34_nl;
  wire LOOPK1_and_156_nl;
  wire LOOPK2_if_1_or_32_nl;
  wire LOOPK1_and_71_nl;
  wire LOOPK2_if_1_or_30_nl;
  wire LOOPK1_and_154_nl;
  wire LOOPK2_if_1_or_28_nl;
  wire LOOPK1_and_69_nl;
  wire LOOPK2_if_1_or_26_nl;
  wire LOOPK1_and_152_nl;
  wire LOOPK2_if_1_or_24_nl;
  wire LOOPK1_and_67_nl;
  wire LOOPK2_if_1_or_22_nl;
  wire LOOPK1_and_150_nl;
  wire LOOPK2_if_1_or_20_nl;
  wire LOOPK1_and_65_nl;
  wire LOOPK2_if_1_or_18_nl;
  wire LOOPK1_and_148_nl;
  wire LOOPK2_if_1_or_16_nl;
  wire LOOPK1_and_81_nl;
  wire LOOPK2_if_1_or_50_nl;
  wire LOOPK1_and_63_nl;
  wire LOOPK2_if_1_or_14_nl;
  wire LOOPK1_and_146_nl;
  wire LOOPK2_if_1_or_12_nl;
  wire LOOPK1_and_61_nl;
  wire LOOPK2_if_1_or_10_nl;
  wire LOOPK1_and_144_nl;
  wire LOOPK2_if_1_or_8_nl;
  wire LOOPK1_and_59_nl;
  wire LOOPK2_if_1_or_6_nl;
  wire LOOPK1_and_142_nl;
  wire LOOPK2_if_1_or_4_nl;
  wire LOOPK1_and_57_nl;
  wire LOOPK2_if_1_or_2_nl;
  wire LOOPK1_and_140_nl;
  wire LOOPK2_if_1_or_nl;
  wire LOOPK1_and_56_nl;
  wire LOOPK2_if_1_or_1_nl;
  wire LOOPK1_and_141_nl;
  wire LOOPK2_if_1_or_3_nl;
  wire LOOPK1_and_164_nl;
  wire LOOPK2_if_1_or_48_nl;
  wire LOOPK1_and_58_nl;
  wire LOOPK2_if_1_or_5_nl;
  wire LOOPK1_and_143_nl;
  wire LOOPK2_if_1_or_7_nl;
  wire LOOPK1_and_60_nl;
  wire LOOPK2_if_1_or_9_nl;
  wire LOOPK1_and_145_nl;
  wire LOOPK2_if_1_or_11_nl;
  wire LOOPK1_and_62_nl;
  wire LOOPK2_if_1_or_13_nl;
  wire LOOPK1_and_147_nl;
  wire LOOPK2_if_1_or_15_nl;
  wire LOOPK1_and_64_nl;
  wire LOOPK2_if_1_or_17_nl;
  wire LOOPK1_and_149_nl;
  wire LOOPK2_if_1_or_19_nl;
  wire LOOPK1_and_66_nl;
  wire LOOPK2_if_1_or_21_nl;
  wire LOOPK1_and_151_nl;
  wire LOOPK2_if_1_or_23_nl;
  wire LOOPK1_and_79_nl;
  wire LOOPK2_if_1_or_46_nl;
  wire LOOPK1_and_68_nl;
  wire LOOPK2_if_1_or_25_nl;
  wire LOOPK1_and_153_nl;
  wire LOOPK2_if_1_or_27_nl;
  wire LOOPK1_and_70_nl;
  wire LOOPK2_if_1_or_29_nl;
  wire LOOPK1_and_155_nl;
  wire LOOPK2_if_1_or_31_nl;
  wire LOOPK1_and_72_nl;
  wire LOOPK2_if_1_or_33_nl;
  wire LOOPK1_and_157_nl;
  wire LOOPK2_if_1_or_35_nl;
  wire LOOPK1_and_74_nl;
  wire LOOPK2_if_1_or_37_nl;
  wire LOOPK1_and_159_nl;
  wire LOOPK2_if_1_or_39_nl;
  wire LOOPK1_and_76_nl;
  wire LOOPK2_if_1_or_41_nl;
  wire LOOPK1_and_161_nl;
  wire LOOPK2_if_1_or_43_nl;
  wire LOOPK1_and_162_nl;
  wire LOOPK2_if_1_or_44_nl;
  wire LOOPK1_and_78_nl;
  wire LOOPK2_if_1_or_45_nl;
  wire LOOPK1_and_163_nl;
  wire LOOPK2_if_1_or_47_nl;
  wire LOOPK1_and_80_nl;
  wire LOOPK2_if_1_or_49_nl;
  wire LOOPK1_and_165_nl;
  wire LOOPK2_if_1_or_51_nl;
  wire LOOPK1_and_82_nl;
  wire LOOPK2_if_1_or_53_nl;
  wire LOOPK1_and_167_nl;
  wire LOOPK2_if_1_or_55_nl;
  wire LOOPK1_and_77_nl;
  wire LOOPK2_if_1_or_42_nl;
  wire LOOPK1_and_160_nl;
  wire LOOPK2_if_1_or_40_nl;
  wire LOOPK1_and_75_nl;
  wire LOOPK2_if_1_or_38_nl;
  wire LOOPK1_and_158_nl;
  wire LOOPK2_if_1_or_36_nl;
  wire avg_not_nl;
  wire LOOPK1_if_LOOPK1_if_and_nl;
  wire[5:0] LOOPI1_i_LOOPI1_i_LOOPI1_i_mux_nl;
  wire LOOPI1_i_and_1_nl;
  wire[13:0] LOOPK2_mux_1_nl;
  wire[13:0] LOOPL1_acc_nl;
  wire[14:0] nl_LOOPL1_acc_nl;
  wire[7:0] LOOPL1_mul_nl;
  wire[3:0] operator_16_true_1_operator_16_true_1_acc_nl;
  wire[4:0] nl_operator_16_true_1_operator_16_true_1_acc_nl;
  wire operator_16_true_1_and_nl;
  wire signed [7:0] nl_LOOPL1_mul_sgnd;
  wire LOOPK2_not_1_nl;
  wire[17:0] operator_20_true_acc_4_nl;
  wire[18:0] nl_operator_20_true_acc_4_nl;
  wire[17:0] LOOPK2_oif_mul_1_nl;
  wire signed [18:0] nl_LOOPK2_oif_mul_1_nl;
  wire or_nl;
  wire mux_4_nl;
  wire[21:0] operator_20_true_acc_nl;
  wire[22:0] nl_operator_20_true_acc_nl;
  wire[14:0] LOOPK2_acc_1_nl;
  wire[15:0] nl_LOOPK2_acc_1_nl;
  wire[4:0] LOOPK2_k_mux_1_nl;
  wire[4:0] LOOPK1_k_LOOPK1_k_and_nl;
  wire LOOPK2_k_not_2_nl;
  wire[3:0] operator_4_false_mux_1_nl;
  wire operator_4_false_or_1_nl;
  wire operator_6_false_operator_6_false_and_2_nl;
  wire operator_6_false_operator_6_false_and_3_nl;
  wire[4:0] operator_6_false_mux_2_nl;
  wire[5:0] operator_7_false_mux_1_nl;
  wire or_287_nl;
  wire[19:0] LOOPK2_mux_3_nl;
  wire[19:0] LOOPK2_oif_mul_2_nl;
  wire signed [20:0] nl_LOOPK2_oif_mul_2_nl;
  wire[19:0] LOOPK2_mux_4_nl;
  wire operator_7_false_operator_7_false_and_2_nl;
  wire[1:0] operator_7_false_operator_7_false_and_3_nl;
  wire[1:0] operator_7_false_mux_1_nl_1;
  wire not_80_nl;
  wire[3:0] operator_7_false_mux1h_3_nl;
  wire or_288_nl;

  // Interconnect Declarations for Component Instantiations 
  wire  nl_ATTENTION_IP_Attention_Filter_run_run_fsm_inst_LOOPK1_C_0_tr0;
  assign nl_ATTENTION_IP_Attention_Filter_run_run_fsm_inst_LOOPK1_C_0_tr0 = mux_tmp_3
      & (~ (z_out_4[6]));
  ATTENTION_IP_Attention_Filter_run_q_chan1_rsci ATTENTION_IP_Attention_Filter_run_q_chan1_rsci_inst
      (
      .q_chan1_rsc_dat(q_chan1_rsc_dat),
      .q_chan1_rsc_vld(q_chan1_rsc_vld),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy),
      .q_chan1_rsci_oswt(reg_q_chan1_rsci_oswt_cse),
      .q_chan1_rsci_wen_comp(q_chan1_rsci_wen_comp),
      .q_chan1_rsci_idat_mxwt(q_chan1_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Filter_run_k_chan1_rsci ATTENTION_IP_Attention_Filter_run_k_chan1_rsci_inst
      (
      .k_chan1_rsc_dat(k_chan1_rsc_dat),
      .k_chan1_rsc_vld(k_chan1_rsc_vld),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy),
      .k_chan1_rsci_oswt(reg_k_chan1_rsci_oswt_cse),
      .k_chan1_rsci_wen_comp(k_chan1_rsci_wen_comp),
      .k_chan1_rsci_idat_mxwt(k_chan1_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Filter_run_v_chan1_rsci ATTENTION_IP_Attention_Filter_run_v_chan1_rsci_inst
      (
      .v_chan1_rsc_dat(v_chan1_rsc_dat),
      .v_chan1_rsc_vld(v_chan1_rsc_vld),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy),
      .v_chan1_rsci_oswt(reg_v_chan1_rsci_oswt_cse),
      .v_chan1_rsci_wen_comp(v_chan1_rsci_wen_comp),
      .v_chan1_rsci_idat_mxwt(v_chan1_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Filter_run_q_chan2_rsci ATTENTION_IP_Attention_Filter_run_q_chan2_rsci_inst
      (
      .q_chan2_rsc_dat(q_chan2_rsc_dat),
      .q_chan2_rsc_vld(q_chan2_rsc_vld),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy),
      .q_chan2_rsci_oswt(reg_q_chan2_rsci_oswt_cse),
      .q_chan2_rsci_wen_comp(q_chan2_rsci_wen_comp),
      .q_chan2_rsci_idat(q_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_k_chan2_rsci ATTENTION_IP_Attention_Filter_run_k_chan2_rsci_inst
      (
      .k_chan2_rsc_dat(k_chan2_rsc_dat),
      .k_chan2_rsc_vld(k_chan2_rsc_vld),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy),
      .k_chan2_rsci_oswt(reg_k_chan2_rsci_oswt_cse),
      .k_chan2_rsci_wen_comp(k_chan2_rsci_wen_comp),
      .k_chan2_rsci_idat(k_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_v_chan2_rsci ATTENTION_IP_Attention_Filter_run_v_chan2_rsci_inst
      (
      .v_chan2_rsc_dat(v_chan2_rsc_dat),
      .v_chan2_rsc_vld(v_chan2_rsc_vld),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy),
      .v_chan2_rsci_oswt(reg_v_chan2_rsci_oswt_cse),
      .v_chan2_rsci_wen_comp(v_chan2_rsci_wen_comp),
      .v_chan2_rsci_idat(v_chan2_rsci_idat)
    );
  ATTENTION_IP_Attention_Filter_run_staller ATTENTION_IP_Attention_Filter_run_staller_inst
      (
      .run_wen(run_wen),
      .q_chan1_rsci_wen_comp(q_chan1_rsci_wen_comp),
      .k_chan1_rsci_wen_comp(k_chan1_rsci_wen_comp),
      .v_chan1_rsci_wen_comp(v_chan1_rsci_wen_comp),
      .q_chan2_rsci_wen_comp(q_chan2_rsci_wen_comp),
      .k_chan2_rsci_wen_comp(k_chan2_rsci_wen_comp),
      .v_chan2_rsci_wen_comp(v_chan2_rsci_wen_comp)
    );
  ATTENTION_IP_Attention_Filter_run_run_fsm ATTENTION_IP_Attention_Filter_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .LOOPI1_C_0_tr0(and_cse),
      .LOOPK1_C_0_tr0(nl_ATTENTION_IP_Attention_Filter_run_run_fsm_inst_LOOPK1_C_0_tr0),
      .LOOPL1_C_0_tr0(LOOPL1_LOOPL1_if_LOOPL1_if_nor_tmp),
      .LOOPK2_C_3_tr0(LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp),
      .LOOPK3_C_1_tr0(LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt),
      .LOOPJ1_C_4_tr0(LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp),
      .LOOPI2_C_0_tr0(LOOPI2_LOOPI2_if_LOOPI2_if_nor_tmp)
    );
  assign LOOPK2_if_1_or_56_itm = and_50_cse | and_52_cse;
  assign sel_and_1_cse = run_wen & ((fsm_output[4]) | and_50_cse);
  assign sel_and_2_cse = run_wen & (((or_tmp_11 | (z_out_4[6])) & (fsm_output[4]))
      | and_50_cse);
  assign and_cse = ~((LOOPI1_i_1_6_1_sva != (z_out_4[6:1])) | (z_out_4[7]));
  assign LOOPK2_if_1_LOOPK2_if_1_nor_2_cse = ~(LOOPK2_k_sva_rsp_0 | (LOOPK2_k_sva_rsp_1!=5'b00000));
  assign LOOPL1_l_nand_seb = ~((~((fsm_output[12]) | (fsm_output[8]))) & (~((fsm_output[7])
      | (fsm_output[9]))));
  assign LOOPI1_i_LOOPI1_i_LOOPI1_i_nor_cse = ~((fsm_output[9:8]!=2'b00));
  assign or_7_cse = LOOPK2_k_sva_rsp_0 | (LOOPK2_k_sva_rsp_1!=5'b00000);
  assign LOOPK1_if_equal_tmp = LOOPK2_k_sva_rsp_1 == (z_out_4[5:1]);
  assign LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp = ~((({LOOPK2_k_sva_rsp_0 , LOOPK2_k_sva_rsp_1})
      != (z_out_4[5:0])) | (z_out_4[6]));
  assign LOOPK1_and_stg_3_1_sva_1 = LOOPK1_and_stg_2_1_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_2_sva_1 = LOOPK1_and_stg_2_2_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_3_sva_1 = LOOPK1_and_stg_2_3_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_4_sva_1 = LOOPK1_and_stg_2_4_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_5_sva_1 = LOOPK1_and_stg_2_5_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_6_sva_1 = LOOPK1_and_stg_2_6_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_7_sva_1 = LOOPK1_and_stg_2_7_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK1_and_stg_3_8_sva_1 = LOOPK1_and_stg_2_0_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK1_and_stg_3_9_sva_1 = LOOPK1_and_stg_2_1_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK1_and_stg_3_10_sva_1 = LOOPK1_and_stg_2_2_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK1_and_stg_3_11_sva_1 = LOOPK1_and_stg_2_3_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK1_and_stg_2_4_sva_1 = LOOPK1_and_stg_1_0_sva_1 & (LOOPK2_k_sva_rsp_1[2]);
  assign LOOPK1_and_stg_2_5_sva_1 = LOOPK1_and_stg_1_1_sva_1 & (LOOPK2_k_sva_rsp_1[2]);
  assign LOOPK1_and_stg_2_6_sva_1 = LOOPK1_and_stg_1_2_sva_1 & (LOOPK2_k_sva_rsp_1[2]);
  assign LOOPK1_and_stg_2_7_sva_1 = LOOPK1_and_stg_1_3_sva_1 & (LOOPK2_k_sva_rsp_1[2]);
  assign LOOPK1_and_stg_2_0_sva_1 = LOOPK1_and_stg_1_0_sva_1 & (~ (LOOPK2_k_sva_rsp_1[2]));
  assign LOOPK1_and_stg_2_1_sva_1 = LOOPK1_and_stg_1_1_sva_1 & (~ (LOOPK2_k_sva_rsp_1[2]));
  assign LOOPK1_and_stg_2_2_sva_1 = LOOPK1_and_stg_1_2_sva_1 & (~ (LOOPK2_k_sva_rsp_1[2]));
  assign LOOPK1_and_stg_2_3_sva_1 = LOOPK1_and_stg_1_3_sva_1 & (~ (LOOPK2_k_sva_rsp_1[2]));
  assign LOOPK1_and_stg_1_0_sva_1 = ~((LOOPK2_k_sva_rsp_1[1:0]!=2'b00));
  assign LOOPK1_and_stg_1_1_sva_1 = (LOOPK2_k_sva_rsp_1[1:0]==2'b01);
  assign LOOPK1_and_stg_1_2_sva_1 = (LOOPK2_k_sva_rsp_1[1:0]==2'b10);
  assign LOOPK1_and_stg_1_3_sva_1 = (LOOPK2_k_sva_rsp_1[1:0]==2'b11);
  assign LOOPK1_not_127 = ~(LOOPK1_and_stg_3_11_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_129 = ~(LOOPK1_and_stg_3_1_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_131 = ~(LOOPK1_and_stg_3_10_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_133 = ~(LOOPK1_and_stg_3_2_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_135 = ~(LOOPK1_and_stg_3_9_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_137 = ~(LOOPK1_and_stg_3_3_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_139 = ~(LOOPK1_and_stg_3_8_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_141 = ~(LOOPK1_and_stg_3_4_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_143 = ~(LOOPK1_and_stg_3_7_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_145 = ~(LOOPK1_and_stg_3_5_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_147 = ~(LOOPK1_and_stg_3_6_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_149 = ~(LOOPK1_and_stg_3_6_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_151 = ~(LOOPK1_and_stg_3_5_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_153 = ~(LOOPK1_and_stg_3_7_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_155 = ~(LOOPK1_and_stg_3_4_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_157 = ~(LOOPK1_and_stg_3_8_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_159 = ~(LOOPK1_and_stg_3_3_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_161 = ~(LOOPK1_and_stg_3_9_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_163 = ~(LOOPK1_and_stg_3_2_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_165 = ~(LOOPK1_and_stg_3_10_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_167 = ~(LOOPK1_and_stg_3_1_sva_1 & (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK1_not_169 = ~(LOOPK1_and_stg_3_11_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4])));
  assign LOOPK1_not_171 = ~(LOOPK1_and_stg_2_0_sva_1 & (LOOPK2_k_sva_rsp_1[4:3]==2'b10));
  assign LOOPK1_not_173 = ~(LOOPK1_and_stg_2_4_sva_1 & (LOOPK2_k_sva_rsp_1[4:3]==2'b01));
  assign LOOPK1_not_175 = ~(LOOPK1_and_stg_2_7_sva_1 & (LOOPK2_k_sva_rsp_1[4:3]==2'b01));
  assign LOOPK1_not_177 = ~(LOOPK1_and_stg_2_5_sva_1 & (LOOPK2_k_sva_rsp_1[4:3]==2'b01));
  assign LOOPK1_not_179 = ~(LOOPK1_and_stg_2_6_sva_1 & (LOOPK2_k_sva_rsp_1[4:3]==2'b01));
  assign operator_16_true_slc_q_channel_data_16_15_0_tmp_sva_1 = MUX_v_16_64_2((q_channel_data_sva[15:0]),
      (q_channel_data_sva[31:16]), (q_channel_data_sva[47:32]), (q_channel_data_sva[63:48]),
      (q_channel_data_sva[79:64]), (q_channel_data_sva[95:80]), (q_channel_data_sva[111:96]),
      (q_channel_data_sva[127:112]), (q_channel_data_sva[143:128]), (q_channel_data_sva[159:144]),
      (q_channel_data_sva[175:160]), (q_channel_data_sva[191:176]), (q_channel_data_sva[207:192]),
      (q_channel_data_sva[223:208]), (q_channel_data_sva[239:224]), (q_channel_data_sva[255:240]),
      (q_channel_data_sva[271:256]), (q_channel_data_sva[287:272]), (q_channel_data_sva[303:288]),
      (q_channel_data_sva[319:304]), (q_channel_data_sva[335:320]), (q_channel_data_sva[351:336]),
      (q_channel_data_sva[367:352]), (q_channel_data_sva[383:368]), (q_channel_data_sva[399:384]),
      (q_channel_data_sva[415:400]), (q_channel_data_sva[431:416]), (q_channel_data_sva[447:432]),
      (q_channel_data_sva[463:448]), (q_channel_data_sva[479:464]), (q_channel_data_sva[495:480]),
      (q_channel_data_sva[511:496]), (q_channel_data_sva[527:512]), (q_channel_data_sva[543:528]),
      (q_channel_data_sva[559:544]), (q_channel_data_sva[575:560]), (q_channel_data_sva[591:576]),
      (q_channel_data_sva[607:592]), (q_channel_data_sva[623:608]), (q_channel_data_sva[639:624]),
      (q_channel_data_sva[655:640]), (q_channel_data_sva[671:656]), (q_channel_data_sva[687:672]),
      (q_channel_data_sva[703:688]), (q_channel_data_sva[719:704]), (q_channel_data_sva[735:720]),
      (q_channel_data_sva[751:736]), (q_channel_data_sva[767:752]), (q_channel_data_sva[783:768]),
      (q_channel_data_sva[799:784]), (q_channel_data_sva[815:800]), (q_channel_data_sva[831:816]),
      (q_channel_data_sva[847:832]), (q_channel_data_sva[863:848]), (q_channel_data_sva[879:864]),
      (q_channel_data_sva[895:880]), (q_channel_data_sva[911:896]), (q_channel_data_sva[927:912]),
      (q_channel_data_sva[943:928]), (q_channel_data_sva[959:944]), (q_channel_data_sva[975:960]),
      (q_channel_data_sva[991:976]), (q_channel_data_sva[1007:992]), (q_channel_data_sva[1023:1008]),
      LOOPL1_l_sva_5_0);
  assign operator_16_true_1_slc_k_channel_data_16_15_0_tmp_sva_1 = MUX_v_16_64_2((k_channel_data_sva[15:0]),
      (k_channel_data_sva[31:16]), (k_channel_data_sva[47:32]), (k_channel_data_sva[63:48]),
      (k_channel_data_sva[79:64]), (k_channel_data_sva[95:80]), (k_channel_data_sva[111:96]),
      (k_channel_data_sva[127:112]), (k_channel_data_sva[143:128]), (k_channel_data_sva[159:144]),
      (k_channel_data_sva[175:160]), (k_channel_data_sva[191:176]), (k_channel_data_sva[207:192]),
      (k_channel_data_sva[223:208]), (k_channel_data_sva[239:224]), (k_channel_data_sva[255:240]),
      (k_channel_data_sva[271:256]), (k_channel_data_sva[287:272]), (k_channel_data_sva[303:288]),
      (k_channel_data_sva[319:304]), (k_channel_data_sva[335:320]), (k_channel_data_sva[351:336]),
      (k_channel_data_sva[367:352]), (k_channel_data_sva[383:368]), (k_channel_data_sva[399:384]),
      (k_channel_data_sva[415:400]), (k_channel_data_sva[431:416]), (k_channel_data_sva[447:432]),
      (k_channel_data_sva[463:448]), (k_channel_data_sva[479:464]), (k_channel_data_sva[495:480]),
      (k_channel_data_sva[511:496]), (k_channel_data_sva[527:512]), (k_channel_data_sva[543:528]),
      (k_channel_data_sva[559:544]), (k_channel_data_sva[575:560]), (k_channel_data_sva[591:576]),
      (k_channel_data_sva[607:592]), (k_channel_data_sva[623:608]), (k_channel_data_sva[639:624]),
      (k_channel_data_sva[655:640]), (k_channel_data_sva[671:656]), (k_channel_data_sva[687:672]),
      (k_channel_data_sva[703:688]), (k_channel_data_sva[719:704]), (k_channel_data_sva[735:720]),
      (k_channel_data_sva[751:736]), (k_channel_data_sva[767:752]), (k_channel_data_sva[783:768]),
      (k_channel_data_sva[799:784]), (k_channel_data_sva[815:800]), (k_channel_data_sva[831:816]),
      (k_channel_data_sva[847:832]), (k_channel_data_sva[863:848]), (k_channel_data_sva[879:864]),
      (k_channel_data_sva[895:880]), (k_channel_data_sva[911:896]), (k_channel_data_sva[927:912]),
      (k_channel_data_sva[943:928]), (k_channel_data_sva[959:944]), (k_channel_data_sva[975:960]),
      (k_channel_data_sva[991:976]), (k_channel_data_sva[1007:992]), (k_channel_data_sva[1023:1008]),
      LOOPL1_l_sva_5_0);
  assign LOOPK2_if_1_and_stg_4_23_sva_1 = LOOPK1_and_stg_3_7_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_22_sva_1 = LOOPK1_and_stg_3_6_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_21_sva_1 = LOOPK1_and_stg_3_5_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_20_sva_1 = LOOPK1_and_stg_3_4_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_19_sva_1 = LOOPK1_and_stg_3_3_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_18_sva_1 = LOOPK1_and_stg_3_2_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_17_sva_1 = LOOPK1_and_stg_3_1_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_16_sva_1 = LOOPK2_if_1_and_stg_3_0_sva_1 & (LOOPK2_k_sva_rsp_1[4]);
  assign LOOPK2_if_1_and_stg_4_15_sva_1 = LOOPK2_if_1_and_stg_3_15_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_14_sva_1 = LOOPK2_if_1_and_stg_3_14_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_13_sva_1 = LOOPK2_if_1_and_stg_3_13_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_12_sva_1 = LOOPK2_if_1_and_stg_3_12_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_11_sva_1 = LOOPK1_and_stg_3_11_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_10_sva_1 = LOOPK1_and_stg_3_10_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_9_sva_1 = LOOPK1_and_stg_3_9_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_8_sva_1 = LOOPK1_and_stg_3_8_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_7_sva_1 = LOOPK1_and_stg_3_7_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_6_sva_1 = LOOPK1_and_stg_3_6_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_5_sva_1 = LOOPK1_and_stg_3_5_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_4_sva_1 = LOOPK1_and_stg_3_4_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_3_sva_1 = LOOPK1_and_stg_3_3_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_2_sva_1 = LOOPK1_and_stg_3_2_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_4_1_sva_1 = LOOPK1_and_stg_3_1_sva_1 & (~ (LOOPK2_k_sva_rsp_1[4]));
  assign LOOPK2_if_1_and_stg_3_0_sva_1 = LOOPK1_and_stg_2_0_sva_1 & (~ (LOOPK2_k_sva_rsp_1[3]));
  assign LOOPK2_if_1_and_stg_3_15_sva_1 = LOOPK1_and_stg_2_7_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK2_if_1_and_stg_3_14_sva_1 = LOOPK1_and_stg_2_6_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK2_if_1_and_stg_3_13_sva_1 = LOOPK1_and_stg_2_5_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPK2_if_1_and_stg_3_12_sva_1 = LOOPK1_and_stg_2_4_sva_1 & (LOOPK2_k_sva_rsp_1[3]);
  assign LOOPI2_LOOPI2_if_LOOPI2_if_nor_tmp = ~((LOOPI2_i_sva != (z_out_4[3:0]))
      | (z_out_4[4]));
  assign LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp = ~((LOOPI1_i_1_6_1_sva != (z_out_4[5:0]))
      | (z_out_4[6]));
  assign LOOPK3_if_1_mux_tmp = MUX_s_1_56_2(1'b1, sel_1_lpi_3, sel_2_lpi_3, sel_3_lpi_3,
      sel_4_lpi_3, sel_5_lpi_3, sel_6_lpi_3, sel_7_lpi_3, sel_8_lpi_3, sel_9_lpi_3,
      sel_10_lpi_3, sel_11_lpi_3, sel_12_lpi_3, sel_13_lpi_3, sel_14_lpi_3, sel_15_lpi_3,
      sel_16_lpi_3, sel_17_lpi_3, sel_18_lpi_3, sel_19_lpi_3, sel_20_lpi_3, sel_21_lpi_3,
      sel_22_lpi_3, sel_23_lpi_3, sel_24_lpi_3, sel_25_lpi_3, sel_26_lpi_3, sel_27_lpi_3,
      sel_28_lpi_3, sel_29_lpi_3, sel_30_lpi_3, sel_31_lpi_3, sel_32_lpi_3, sel_33_lpi_3,
      sel_34_lpi_3, sel_35_lpi_3, sel_36_lpi_3, sel_37_lpi_3, sel_38_lpi_3, sel_39_lpi_3,
      sel_40_lpi_3, sel_41_lpi_3, sel_42_lpi_3, sel_43_lpi_3, sel_44_lpi_3, sel_45_lpi_3,
      sel_46_lpi_3, sel_47_lpi_3, sel_48_lpi_3, sel_49_lpi_3, sel_50_lpi_3, sel_51_lpi_3,
      sel_52_lpi_3, sel_53_lpi_3, sel_54_lpi_3, sel_55_lpi_3, {LOOPK2_k_sva_rsp_0
      , LOOPK2_k_sva_rsp_1});
  assign LOOPL1_LOOPL1_if_LOOPL1_if_nor_tmp = ~((({LOOPL1_l_sva_6 , LOOPL1_l_sva_5_0})
      != (z_out_4[6:0])) | (z_out_4[7]));
  assign LOOPK1_if_unequal_tmp = LOOPK2_k_sva_rsp_1 != (z_out_4[5:1]);
  assign or_tmp_11 = LOOPK1_if_unequal_tmp | (z_out_4[0]);
  assign or_nl = (z_out_4[0]) | (~ LOOPK1_if_unequal_tmp);
  assign mux_tmp_3 = MUX_s_1_2_2((~ or_tmp_11), or_nl, LOOPK1_if_equal_tmp);
  assign nl_operator_20_true_acc_nl = conv_s2u_21_22({operator_20_true_acc_3_itm_21_2
      , (avg_sva[0])}) + conv_s2u_20_22(z_out_3[20:1]);
  assign operator_20_true_acc_nl = nl_operator_20_true_acc_nl[21:0];
  assign mux_4_nl = MUX_s_1_2_2(LOOPK2_if_1_LOOPK2_if_1_nor_2_cse, or_7_cse, readslicef_22_1_21(operator_20_true_acc_nl));
  assign and_50_cse = (mux_4_nl | LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt) & (fsm_output[9]);
  assign and_52_cse = LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp & (fsm_output[10]);
  assign and_65_cse = and_cse & (fsm_output[1]);
  assign or_tmp_198 = (~((fsm_output[8:6]!=3'b000))) & (~((fsm_output[4]) | (fsm_output[5])
      | (fsm_output[10])));
  assign LOOPI1_i_1_6_1_sva_mx0c1 = (fsm_output[0]) | (fsm_output[15]) | and_65_cse;
  assign sel_1_lpi_3_mx0c0 = ((~ mux_tmp_3) | (z_out_4[6])) & (fsm_output[4]);
  assign LOOPK2_k_sva_mx0c1 = (fsm_output[11]) | (fsm_output[5]);
  assign LOOPK2_k_sva_mx0c2 = (fsm_output[13]) | (fsm_output[10]);
  assign nl_LOOPK2_acc_1_nl = conv_s2u_14_15(max_sva) - conv_s2u_14_15(LOOPK2_mux_106_itm);
  assign LOOPK2_acc_1_nl = nl_LOOPK2_acc_1_nl[14:0];
  assign LOOPK2_mux_106_itm_mx0c2 = (~ (readslicef_15_1_14(LOOPK2_acc_1_nl))) & (fsm_output[8]);
  assign or_282_itm = (fsm_output[10]) | (fsm_output[14]) | (fsm_output[4]) | (fsm_output[12]);
  assign LOOPK2_k_and_ssc = run_wen & ((fsm_output[4:3]!=2'b00) | LOOPK2_k_sva_mx0c1
      | LOOPK2_k_sva_mx0c2);
  always @(posedge clk) begin
    if ( run_wen & LOOPK2_if_1_or_56_itm ) begin
      k_chan2_rsci_idat <= MUX_v_1024_2_2(1024'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000,
          k_channel_data_sva, LOOPK2_if_1_not_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[12]) & LOOPK3_if_1_mux_tmp ) begin
      v_chan2_rsci_idat <= v_chan1_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[2]) ) begin
      q_chan2_rsci_idat <= q_chan1_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & ((fsm_output[1]) | (fsm_output[14]) | LOOPI1_i_1_6_1_sva_mx0c1)
        ) begin
      LOOPI1_i_1_6_1_sva <= MUX_v_6_2_2(6'b000000, z_out_2, LOOPI1_i_not_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_q_chan1_rsci_oswt_cse <= 1'b0;
      reg_k_chan1_rsci_oswt_cse <= 1'b0;
      reg_v_chan1_rsci_oswt_cse <= 1'b0;
      reg_q_chan2_rsci_oswt_cse <= 1'b0;
      reg_k_chan2_rsci_oswt_cse <= 1'b0;
      reg_v_chan2_rsci_oswt_cse <= 1'b0;
      LOOPL1_l_sva_6 <= 1'b0;
    end
    else if ( rst ) begin
      reg_q_chan1_rsci_oswt_cse <= 1'b0;
      reg_k_chan1_rsci_oswt_cse <= 1'b0;
      reg_v_chan1_rsci_oswt_cse <= 1'b0;
      reg_q_chan2_rsci_oswt_cse <= 1'b0;
      reg_k_chan2_rsci_oswt_cse <= 1'b0;
      reg_v_chan2_rsci_oswt_cse <= 1'b0;
      LOOPL1_l_sva_6 <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_q_chan1_rsci_oswt_cse <= ((~ LOOPI2_LOOPI2_if_LOOPI2_if_nor_tmp) & (fsm_output[15]))
          | and_65_cse | ((~ LOOPJ1_LOOPJ1_if_1_LOOPJ1_if_1_nor_tmp) & (fsm_output[14]));
      reg_k_chan1_rsci_oswt_cse <= (fsm_output[5]) | ((~ LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp)
          & (fsm_output[10]));
      reg_v_chan1_rsci_oswt_cse <= (fsm_output[11]) | ((~ LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt)
          & (fsm_output[13]));
      reg_q_chan2_rsci_oswt_cse <= fsm_output[2];
      reg_k_chan2_rsci_oswt_cse <= LOOPK2_if_1_or_56_itm;
      reg_v_chan2_rsci_oswt_cse <= LOOPK3_if_1_mux_tmp & (fsm_output[12]);
      LOOPL1_l_sva_6 <= (z_out_1[6]) & LOOPL1_l_nand_seb;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (sel_1_lpi_3_mx0c0 | (fsm_output[5]) | and_50_cse) ) begin
      sel_1_lpi_3 <= ~(sel_mux_nl | sel_1_lpi_3_mx0c0);
    end
  end
  always @(posedge clk) begin
    if ( sel_and_1_cse ) begin
      sel_10_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_73_nl, LOOPK2_if_1_or_34_nl, and_50_cse);
      sel_12_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_71_nl, LOOPK2_if_1_or_30_nl, and_50_cse);
      sel_14_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_69_nl, LOOPK2_if_1_or_26_nl, and_50_cse);
      sel_16_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_67_nl, LOOPK2_if_1_or_22_nl, and_50_cse);
      sel_18_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_65_nl, LOOPK2_if_1_or_18_nl, and_50_cse);
      sel_2_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_81_nl, LOOPK2_if_1_or_50_nl, and_50_cse);
      sel_20_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_63_nl, LOOPK2_if_1_or_14_nl, and_50_cse);
      sel_22_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_61_nl, LOOPK2_if_1_or_10_nl, and_50_cse);
      sel_24_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_59_nl, LOOPK2_if_1_or_6_nl, and_50_cse);
      sel_26_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_57_nl, LOOPK2_if_1_or_2_nl, and_50_cse);
      sel_28_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_56_nl, LOOPK2_if_1_or_1_nl, and_50_cse);
      sel_30_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_58_nl, LOOPK2_if_1_or_5_nl, and_50_cse);
      sel_32_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_60_nl, LOOPK2_if_1_or_9_nl, and_50_cse);
      sel_34_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_62_nl, LOOPK2_if_1_or_13_nl, and_50_cse);
      sel_36_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_64_nl, LOOPK2_if_1_or_17_nl, and_50_cse);
      sel_38_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_66_nl, LOOPK2_if_1_or_21_nl, and_50_cse);
      sel_4_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_79_nl, LOOPK2_if_1_or_46_nl, and_50_cse);
      sel_40_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_68_nl, LOOPK2_if_1_or_25_nl, and_50_cse);
      sel_42_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_70_nl, LOOPK2_if_1_or_29_nl, and_50_cse);
      sel_44_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_72_nl, LOOPK2_if_1_or_33_nl, and_50_cse);
      sel_46_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_74_nl, LOOPK2_if_1_or_37_nl, and_50_cse);
      sel_48_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_76_nl, LOOPK2_if_1_or_41_nl, and_50_cse);
      sel_50_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_78_nl, LOOPK2_if_1_or_45_nl, and_50_cse);
      sel_52_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_80_nl, LOOPK2_if_1_or_49_nl, and_50_cse);
      sel_54_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_82_nl, LOOPK2_if_1_or_53_nl, and_50_cse);
      sel_6_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_77_nl, LOOPK2_if_1_or_42_nl, and_50_cse);
      sel_8_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_75_nl, LOOPK2_if_1_or_38_nl, and_50_cse);
    end
  end
  always @(posedge clk) begin
    if ( sel_and_2_cse ) begin
      sel_11_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_156_nl, LOOPK2_if_1_or_32_nl, and_50_cse);
      sel_13_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_154_nl, LOOPK2_if_1_or_28_nl, and_50_cse);
      sel_15_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_152_nl, LOOPK2_if_1_or_24_nl, and_50_cse);
      sel_17_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_150_nl, LOOPK2_if_1_or_20_nl, and_50_cse);
      sel_19_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_148_nl, LOOPK2_if_1_or_16_nl, and_50_cse);
      sel_21_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_146_nl, LOOPK2_if_1_or_12_nl, and_50_cse);
      sel_23_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_144_nl, LOOPK2_if_1_or_8_nl, and_50_cse);
      sel_25_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_142_nl, LOOPK2_if_1_or_4_nl, and_50_cse);
      sel_27_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_140_nl, LOOPK2_if_1_or_nl, and_50_cse);
      sel_29_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_141_nl, LOOPK2_if_1_or_3_nl, and_50_cse);
      sel_3_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_164_nl, LOOPK2_if_1_or_48_nl, and_50_cse);
      sel_31_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_143_nl, LOOPK2_if_1_or_7_nl, and_50_cse);
      sel_33_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_145_nl, LOOPK2_if_1_or_11_nl, and_50_cse);
      sel_35_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_147_nl, LOOPK2_if_1_or_15_nl, and_50_cse);
      sel_37_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_149_nl, LOOPK2_if_1_or_19_nl, and_50_cse);
      sel_39_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_151_nl, LOOPK2_if_1_or_23_nl, and_50_cse);
      sel_41_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_153_nl, LOOPK2_if_1_or_27_nl, and_50_cse);
      sel_43_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_155_nl, LOOPK2_if_1_or_31_nl, and_50_cse);
      sel_45_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_157_nl, LOOPK2_if_1_or_35_nl, and_50_cse);
      sel_47_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_159_nl, LOOPK2_if_1_or_39_nl, and_50_cse);
      sel_49_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_161_nl, LOOPK2_if_1_or_43_nl, and_50_cse);
      sel_5_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_162_nl, LOOPK2_if_1_or_44_nl, and_50_cse);
      sel_51_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_163_nl, LOOPK2_if_1_or_47_nl, and_50_cse);
      sel_53_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_165_nl, LOOPK2_if_1_or_51_nl, and_50_cse);
      sel_55_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_167_nl, LOOPK2_if_1_or_55_nl, and_50_cse);
      sel_7_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_160_nl, LOOPK2_if_1_or_40_nl, and_50_cse);
      sel_9_lpi_3 <= MUX_s_1_2_2(LOOPK1_and_158_nl, LOOPK2_if_1_or_36_nl, and_50_cse);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & ((fsm_output[1]) | (fsm_output[15])) ) begin
      LOOPI2_i_sva <= MUX_v_4_2_2(4'b0000, z_out, (fsm_output[15]));
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[10:3]==8'b00000000) ) begin
      q_channel_data_sva <= q_chan1_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( (fsm_output[8:4]==5'b00000) & run_wen ) begin
      avg_sva <= MUX_v_20_2_2(20'b00000000000000000000, LOOPK2_acc_2_itm, avg_not_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (or_tmp_198 | (fsm_output[10])) ) begin
      max_sva <= MUX_v_14_2_2(14'b10000000000000, LOOPK2_mux_106_itm, fsm_output[10]);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt <= 1'b0;
    end
    else if ( rst ) begin
      LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt <= 1'b0;
    end
    else if ( run_wen & ((fsm_output[12]) | (fsm_output[7]) | (fsm_output[4])) )
        begin
      LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt <= MUX1HOT_s_1_3_2(LOOPK1_if_LOOPK1_if_and_nl,
          LOOPK2_if_1_LOOPK2_if_1_nor_2_cse, LOOPK3_LOOPK3_if_2_LOOPK3_if_2_nor_tmp,
          {(fsm_output[4]) , (fsm_output[7]) , (fsm_output[12])});
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[8:7]==2'b00) ) begin
      k_channel_data_sva <= k_chan1_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPL1_l_sva_5_0 <= 6'b000000;
    end
    else if ( rst ) begin
      LOOPL1_l_sva_5_0 <= 6'b000000;
    end
    else if ( LOOPI1_i_LOOPI1_i_LOOPI1_i_nor_cse & run_wen ) begin
      LOOPL1_l_sva_5_0 <= MUX_v_6_2_2(6'b000000, LOOPI1_i_LOOPI1_i_LOOPI1_i_mux_nl,
          LOOPL1_l_nand_seb);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & ((fsm_output[7:6]!=2'b00) | LOOPK2_mux_106_itm_mx0c2) ) begin
      LOOPK2_mux_106_itm <= MUX_v_14_2_2(14'b00000000000000, LOOPK2_mux_1_nl, LOOPK2_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & or_7_cse ) begin
      operator_20_true_acc_3_itm_21_2 <= nl_operator_20_true_acc_3_itm_21_2[19:0];
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (fsm_output[8]) ) begin
      LOOPK2_acc_2_itm <= z_out_3[19:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPK2_k_sva_rsp_0 <= 1'b0;
      LOOPK2_k_sva_rsp_1 <= 5'b00000;
    end
    else if ( rst ) begin
      LOOPK2_k_sva_rsp_0 <= 1'b0;
      LOOPK2_k_sva_rsp_1 <= 5'b00000;
    end
    else if ( LOOPK2_k_and_ssc ) begin
      LOOPK2_k_sva_rsp_0 <= (LOOPL1_l_sva_5_0[5]) & (~ LOOPK2_k_sva_mx0c1);
      LOOPK2_k_sva_rsp_1 <= MUX_v_5_2_2(5'b00000, LOOPK2_k_mux_1_nl, LOOPK2_k_not_2_nl);
    end
  end
  assign LOOPK2_if_1_not_nl = ~ and_52_cse;
  assign LOOPI1_i_not_nl = ~ LOOPI1_i_1_6_1_sva_mx0c1;
  assign sel_nand_nl = ~(sel_1_lpi_3 & (~ LOOPK1_2_LOOPK1_if_LOOPK1_if_nor_sxt));
  assign sel_nor_nl = ~(sel_1_lpi_3 | (LOOPK2_if_1_and_stg_4_1_sva_1 & (~ LOOPK2_k_sva_rsp_0)));
  assign sel_mux_nl = MUX_s_1_2_2(sel_nand_nl, sel_nor_nl, and_50_cse);
  assign LOOPK1_and_73_nl = sel_10_lpi_3 & LOOPK1_not_145;
  assign LOOPK2_if_1_or_34_nl = sel_10_lpi_3 | (LOOPK2_if_1_and_stg_4_10_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_71_nl = sel_12_lpi_3 & LOOPK1_not_149;
  assign LOOPK2_if_1_or_30_nl = sel_12_lpi_3 | (LOOPK2_if_1_and_stg_4_12_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_69_nl = sel_14_lpi_3 & LOOPK1_not_153;
  assign LOOPK2_if_1_or_26_nl = sel_14_lpi_3 | (LOOPK2_if_1_and_stg_4_14_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_67_nl = sel_16_lpi_3 & LOOPK1_not_157;
  assign LOOPK2_if_1_or_22_nl = sel_16_lpi_3 | (LOOPK2_if_1_and_stg_4_16_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_65_nl = sel_18_lpi_3 & LOOPK1_not_161;
  assign LOOPK2_if_1_or_18_nl = sel_18_lpi_3 | (LOOPK2_if_1_and_stg_4_18_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_81_nl = sel_2_lpi_3 & LOOPK1_not_129;
  assign LOOPK2_if_1_or_50_nl = sel_2_lpi_3 | (LOOPK2_if_1_and_stg_4_2_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_63_nl = sel_20_lpi_3 & LOOPK1_not_165;
  assign LOOPK2_if_1_or_14_nl = sel_20_lpi_3 | (LOOPK2_if_1_and_stg_4_20_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_61_nl = sel_22_lpi_3 & LOOPK1_not_169;
  assign LOOPK2_if_1_or_10_nl = sel_22_lpi_3 | (LOOPK2_if_1_and_stg_4_22_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_59_nl = sel_24_lpi_3 & LOOPK1_not_173;
  assign LOOPK2_if_1_or_6_nl = sel_24_lpi_3 | (LOOPK1_and_stg_3_8_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_57_nl = sel_26_lpi_3 & LOOPK1_not_177;
  assign LOOPK2_if_1_or_2_nl = sel_26_lpi_3 | (LOOPK1_and_stg_3_10_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_56_nl = sel_28_lpi_3 & LOOPK1_not_179;
  assign LOOPK2_if_1_or_1_nl = sel_28_lpi_3 | (LOOPK2_if_1_and_stg_3_12_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_58_nl = sel_30_lpi_3 & LOOPK1_not_175;
  assign LOOPK2_if_1_or_5_nl = sel_30_lpi_3 | (LOOPK2_if_1_and_stg_3_14_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_60_nl = sel_32_lpi_3 & LOOPK1_not_171;
  assign LOOPK2_if_1_or_9_nl = sel_32_lpi_3 | (LOOPK2_if_1_and_stg_3_0_sva_1 & (~
      (LOOPK2_k_sva_rsp_1[4])) & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_62_nl = sel_34_lpi_3 & LOOPK1_not_167;
  assign LOOPK2_if_1_or_13_nl = sel_34_lpi_3 | (LOOPK2_if_1_and_stg_4_2_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_64_nl = sel_36_lpi_3 & LOOPK1_not_163;
  assign LOOPK2_if_1_or_17_nl = sel_36_lpi_3 | (LOOPK2_if_1_and_stg_4_4_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_66_nl = sel_38_lpi_3 & LOOPK1_not_159;
  assign LOOPK2_if_1_or_21_nl = sel_38_lpi_3 | (LOOPK2_if_1_and_stg_4_6_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_79_nl = sel_4_lpi_3 & LOOPK1_not_133;
  assign LOOPK2_if_1_or_46_nl = sel_4_lpi_3 | (LOOPK2_if_1_and_stg_4_4_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_68_nl = sel_40_lpi_3 & LOOPK1_not_155;
  assign LOOPK2_if_1_or_25_nl = sel_40_lpi_3 | (LOOPK2_if_1_and_stg_4_8_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_70_nl = sel_42_lpi_3 & LOOPK1_not_151;
  assign LOOPK2_if_1_or_29_nl = sel_42_lpi_3 | (LOOPK2_if_1_and_stg_4_10_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_72_nl = sel_44_lpi_3 & LOOPK1_not_147;
  assign LOOPK2_if_1_or_33_nl = sel_44_lpi_3 | (LOOPK2_if_1_and_stg_4_12_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_74_nl = sel_46_lpi_3 & LOOPK1_not_143;
  assign LOOPK2_if_1_or_37_nl = sel_46_lpi_3 | (LOOPK2_if_1_and_stg_4_14_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_76_nl = sel_48_lpi_3 & LOOPK1_not_139;
  assign LOOPK2_if_1_or_41_nl = sel_48_lpi_3 | (LOOPK2_if_1_and_stg_4_16_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_78_nl = sel_50_lpi_3 & LOOPK1_not_135;
  assign LOOPK2_if_1_or_45_nl = sel_50_lpi_3 | (LOOPK2_if_1_and_stg_4_18_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_80_nl = sel_52_lpi_3 & LOOPK1_not_131;
  assign LOOPK2_if_1_or_49_nl = sel_52_lpi_3 | (LOOPK2_if_1_and_stg_4_20_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_82_nl = sel_54_lpi_3 & LOOPK1_not_127;
  assign LOOPK2_if_1_or_53_nl = sel_54_lpi_3 | (LOOPK2_if_1_and_stg_4_22_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_77_nl = sel_6_lpi_3 & LOOPK1_not_137;
  assign LOOPK2_if_1_or_42_nl = sel_6_lpi_3 | (LOOPK2_if_1_and_stg_4_6_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_75_nl = sel_8_lpi_3 & LOOPK1_not_141;
  assign LOOPK2_if_1_or_38_nl = sel_8_lpi_3 | (LOOPK2_if_1_and_stg_4_8_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_156_nl = sel_11_lpi_3 & LOOPK1_not_145;
  assign LOOPK2_if_1_or_32_nl = sel_11_lpi_3 | (LOOPK2_if_1_and_stg_4_11_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_154_nl = sel_13_lpi_3 & LOOPK1_not_149;
  assign LOOPK2_if_1_or_28_nl = sel_13_lpi_3 | (LOOPK2_if_1_and_stg_4_13_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_152_nl = sel_15_lpi_3 & LOOPK1_not_153;
  assign LOOPK2_if_1_or_24_nl = sel_15_lpi_3 | (LOOPK2_if_1_and_stg_4_15_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_150_nl = sel_17_lpi_3 & LOOPK1_not_157;
  assign LOOPK2_if_1_or_20_nl = sel_17_lpi_3 | (LOOPK2_if_1_and_stg_4_17_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_148_nl = sel_19_lpi_3 & LOOPK1_not_161;
  assign LOOPK2_if_1_or_16_nl = sel_19_lpi_3 | (LOOPK2_if_1_and_stg_4_19_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_146_nl = sel_21_lpi_3 & LOOPK1_not_165;
  assign LOOPK2_if_1_or_12_nl = sel_21_lpi_3 | (LOOPK2_if_1_and_stg_4_21_sva_1 &
      (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_144_nl = sel_23_lpi_3 & LOOPK1_not_169;
  assign LOOPK2_if_1_or_8_nl = sel_23_lpi_3 | (LOOPK2_if_1_and_stg_4_23_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_142_nl = sel_25_lpi_3 & LOOPK1_not_173;
  assign LOOPK2_if_1_or_4_nl = sel_25_lpi_3 | (LOOPK1_and_stg_3_9_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_140_nl = sel_27_lpi_3 & LOOPK1_not_177;
  assign LOOPK2_if_1_or_nl = sel_27_lpi_3 | (LOOPK1_and_stg_3_11_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_141_nl = sel_29_lpi_3 & LOOPK1_not_179;
  assign LOOPK2_if_1_or_3_nl = sel_29_lpi_3 | (LOOPK2_if_1_and_stg_3_13_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_164_nl = sel_3_lpi_3 & LOOPK1_not_129;
  assign LOOPK2_if_1_or_48_nl = sel_3_lpi_3 | (LOOPK2_if_1_and_stg_4_3_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_143_nl = sel_31_lpi_3 & LOOPK1_not_175;
  assign LOOPK2_if_1_or_7_nl = sel_31_lpi_3 | (LOOPK2_if_1_and_stg_3_15_sva_1 & (LOOPK2_k_sva_rsp_1[4])
      & (~ LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_145_nl = sel_33_lpi_3 & LOOPK1_not_171;
  assign LOOPK2_if_1_or_11_nl = sel_33_lpi_3 | (LOOPK2_if_1_and_stg_4_1_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_147_nl = sel_35_lpi_3 & LOOPK1_not_167;
  assign LOOPK2_if_1_or_15_nl = sel_35_lpi_3 | (LOOPK2_if_1_and_stg_4_3_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_149_nl = sel_37_lpi_3 & LOOPK1_not_163;
  assign LOOPK2_if_1_or_19_nl = sel_37_lpi_3 | (LOOPK2_if_1_and_stg_4_5_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_151_nl = sel_39_lpi_3 & LOOPK1_not_159;
  assign LOOPK2_if_1_or_23_nl = sel_39_lpi_3 | (LOOPK2_if_1_and_stg_4_7_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_153_nl = sel_41_lpi_3 & LOOPK1_not_155;
  assign LOOPK2_if_1_or_27_nl = sel_41_lpi_3 | (LOOPK2_if_1_and_stg_4_9_sva_1 & LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_155_nl = sel_43_lpi_3 & LOOPK1_not_151;
  assign LOOPK2_if_1_or_31_nl = sel_43_lpi_3 | (LOOPK2_if_1_and_stg_4_11_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_157_nl = sel_45_lpi_3 & LOOPK1_not_147;
  assign LOOPK2_if_1_or_35_nl = sel_45_lpi_3 | (LOOPK2_if_1_and_stg_4_13_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_159_nl = sel_47_lpi_3 & LOOPK1_not_143;
  assign LOOPK2_if_1_or_39_nl = sel_47_lpi_3 | (LOOPK2_if_1_and_stg_4_15_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_161_nl = sel_49_lpi_3 & LOOPK1_not_139;
  assign LOOPK2_if_1_or_43_nl = sel_49_lpi_3 | (LOOPK2_if_1_and_stg_4_17_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_162_nl = sel_5_lpi_3 & LOOPK1_not_133;
  assign LOOPK2_if_1_or_44_nl = sel_5_lpi_3 | (LOOPK2_if_1_and_stg_4_5_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_163_nl = sel_51_lpi_3 & LOOPK1_not_135;
  assign LOOPK2_if_1_or_47_nl = sel_51_lpi_3 | (LOOPK2_if_1_and_stg_4_19_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_165_nl = sel_53_lpi_3 & LOOPK1_not_131;
  assign LOOPK2_if_1_or_51_nl = sel_53_lpi_3 | (LOOPK2_if_1_and_stg_4_21_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_167_nl = sel_55_lpi_3 & LOOPK1_not_127;
  assign LOOPK2_if_1_or_55_nl = sel_55_lpi_3 | (LOOPK2_if_1_and_stg_4_23_sva_1 &
      LOOPK2_k_sva_rsp_0);
  assign LOOPK1_and_160_nl = sel_7_lpi_3 & LOOPK1_not_137;
  assign LOOPK2_if_1_or_40_nl = sel_7_lpi_3 | (LOOPK2_if_1_and_stg_4_7_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign LOOPK1_and_158_nl = sel_9_lpi_3 & LOOPK1_not_141;
  assign LOOPK2_if_1_or_36_nl = sel_9_lpi_3 | (LOOPK2_if_1_and_stg_4_9_sva_1 & (~
      LOOPK2_k_sva_rsp_0));
  assign avg_not_nl = ~ or_tmp_198;
  assign LOOPK1_if_LOOPK1_if_and_nl = (~((~ LOOPK1_if_equal_tmp) | (z_out_4[6])))
      & (z_out_4[0]);
  assign LOOPI1_i_and_1_nl = LOOPI1_i_LOOPI1_i_LOOPI1_i_nor_cse & ((LOOPL1_LOOPL1_if_LOOPL1_if_nor_tmp
      & (fsm_output[7])) | (fsm_output[12]) | (fsm_output[8]) | (fsm_output[9]));
  assign LOOPI1_i_LOOPI1_i_LOOPI1_i_mux_nl = MUX_v_6_2_2((z_out_1[5:0]), z_out_2,
      LOOPI1_i_and_1_nl);
  assign operator_16_true_1_and_nl = (operator_16_true_1_slc_k_channel_data_16_15_0_tmp_sva_1[15])
      & ((operator_16_true_1_slc_k_channel_data_16_15_0_tmp_sva_1[11:0]!=12'b000000000000));
  assign nl_operator_16_true_1_operator_16_true_1_acc_nl = (operator_16_true_1_slc_k_channel_data_16_15_0_tmp_sva_1[15:12])
      + conv_u2s_1_4(operator_16_true_1_and_nl);
  assign operator_16_true_1_operator_16_true_1_acc_nl = nl_operator_16_true_1_operator_16_true_1_acc_nl[3:0];
  assign nl_LOOPL1_mul_sgnd = $signed((z_out)) * $signed(operator_16_true_1_operator_16_true_1_acc_nl);
  assign LOOPL1_mul_nl = $unsigned(nl_LOOPL1_mul_sgnd);
  assign nl_LOOPL1_acc_nl = LOOPK2_mux_106_itm + conv_s2s_8_14(LOOPL1_mul_nl);
  assign LOOPL1_acc_nl = nl_LOOPL1_acc_nl[13:0];
  assign LOOPK2_mux_1_nl = MUX_v_14_2_2(LOOPL1_acc_nl, max_sva, LOOPK2_mux_106_itm_mx0c2);
  assign LOOPK2_not_1_nl = ~ (fsm_output[6]);
  assign nl_LOOPK2_oif_mul_1_nl = $signed(conv_u2s_6_7({LOOPK2_k_sva_rsp_0 , LOOPK2_k_sva_rsp_1}))
      * $signed((LOOPK2_mux_106_itm[11:0]));
  assign LOOPK2_oif_mul_1_nl = nl_LOOPK2_oif_mul_1_nl[17:0];
  assign nl_operator_20_true_acc_4_nl =  -LOOPK2_oif_mul_1_nl;
  assign operator_20_true_acc_4_nl = nl_operator_20_true_acc_4_nl[17:0];
  assign nl_operator_20_true_acc_3_itm_21_2  = conv_s2u_19_20(avg_sva[19:1]) + conv_s2u_18_20(operator_20_true_acc_4_nl);
  assign LOOPK1_k_LOOPK1_k_and_nl = MUX_v_5_2_2(5'b00000, (z_out_1[4:0]), (fsm_output[4]));
  assign LOOPK2_k_mux_1_nl = MUX_v_5_2_2(LOOPK1_k_LOOPK1_k_and_nl, (LOOPL1_l_sva_5_0[4:0]),
      LOOPK2_k_sva_mx0c2);
  assign LOOPK2_k_not_2_nl = ~ LOOPK2_k_sva_mx0c1;
  assign operator_4_false_mux_1_nl = MUX_v_4_2_2(LOOPI2_i_sva, (operator_16_true_slc_q_channel_data_16_15_0_tmp_sva_1[15:12]),
      fsm_output[7]);
  assign operator_4_false_or_1_nl = ((operator_16_true_slc_q_channel_data_16_15_0_tmp_sva_1[15])
      & ((operator_16_true_slc_q_channel_data_16_15_0_tmp_sva_1[11:0]!=12'b000000000000)))
      | (fsm_output[15]);
  assign nl_z_out = operator_4_false_mux_1_nl + conv_u2u_1_4(operator_4_false_or_1_nl);
  assign z_out = nl_z_out[3:0];
  assign operator_6_false_operator_6_false_and_2_nl = LOOPL1_l_sva_6 & (fsm_output[7]);
  assign operator_6_false_operator_6_false_and_3_nl = (LOOPL1_l_sva_5_0[5]) & (fsm_output[7]);
  assign operator_6_false_mux_2_nl = MUX_v_5_2_2(LOOPK2_k_sva_rsp_1, (LOOPL1_l_sva_5_0[4:0]),
      fsm_output[7]);
  assign nl_z_out_1 = ({operator_6_false_operator_6_false_and_2_nl , operator_6_false_operator_6_false_and_3_nl
      , operator_6_false_mux_2_nl}) + 7'b0000001;
  assign z_out_1 = nl_z_out_1[6:0];
  assign or_287_nl = (fsm_output[7]) | (fsm_output[12]);
  assign operator_7_false_mux_1_nl = MUX_v_6_2_2(LOOPI1_i_1_6_1_sva, ({LOOPK2_k_sva_rsp_0
      , LOOPK2_k_sva_rsp_1}), or_287_nl);
  assign nl_z_out_2 = operator_7_false_mux_1_nl + 6'b000001;
  assign z_out_2 = nl_z_out_2[5:0];
  assign nl_LOOPK2_oif_mul_2_nl = $signed(max_sva) * $signed(conv_u2s_6_7({LOOPK2_k_sva_rsp_0
      , LOOPK2_k_sva_rsp_1}));
  assign LOOPK2_oif_mul_2_nl = nl_LOOPK2_oif_mul_2_nl[19:0];
  assign LOOPK2_mux_3_nl = MUX_v_20_2_2(avg_sva, LOOPK2_oif_mul_2_nl, fsm_output[9]);
  assign LOOPK2_mux_4_nl = MUX_v_20_2_2(({{6{LOOPK2_mux_106_itm[13]}}, LOOPK2_mux_106_itm}),
      avg_sva, fsm_output[9]);
  assign nl_z_out_3 = conv_s2u_20_21(LOOPK2_mux_3_nl) + conv_s2u_20_21(LOOPK2_mux_4_nl);
  assign z_out_3 = nl_z_out_3[20:0];
  assign operator_7_false_operator_7_false_and_2_nl = (dim[6]) & (~(or_282_itm |
      (fsm_output[15])));
  assign operator_7_false_mux_1_nl_1 = MUX_v_2_2_2((dim[5:4]), (length[5:4]), or_282_itm);
  assign not_80_nl = ~ (fsm_output[15]);
  assign operator_7_false_operator_7_false_and_3_nl = MUX_v_2_2_2(2'b00, operator_7_false_mux_1_nl_1,
      not_80_nl);
  assign or_288_nl = (fsm_output[7]) | (fsm_output[1]);
  assign operator_7_false_mux1h_3_nl = MUX1HOT_v_4_3_2((dim[3:0]), (length[3:0]),
      head, {or_288_nl , or_282_itm , (fsm_output[15])});
  assign nl_z_out_4 = conv_u2u_7_8({operator_7_false_operator_7_false_and_2_nl ,
      operator_7_false_operator_7_false_and_3_nl , operator_7_false_mux1h_3_nl})
      + 8'b11111111;
  assign z_out_4 = nl_z_out_4[7:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_56_2;
    input  input_0;
    input  input_1;
    input  input_2;
    input  input_3;
    input  input_4;
    input  input_5;
    input  input_6;
    input  input_7;
    input  input_8;
    input  input_9;
    input  input_10;
    input  input_11;
    input  input_12;
    input  input_13;
    input  input_14;
    input  input_15;
    input  input_16;
    input  input_17;
    input  input_18;
    input  input_19;
    input  input_20;
    input  input_21;
    input  input_22;
    input  input_23;
    input  input_24;
    input  input_25;
    input  input_26;
    input  input_27;
    input  input_28;
    input  input_29;
    input  input_30;
    input  input_31;
    input  input_32;
    input  input_33;
    input  input_34;
    input  input_35;
    input  input_36;
    input  input_37;
    input  input_38;
    input  input_39;
    input  input_40;
    input  input_41;
    input  input_42;
    input  input_43;
    input  input_44;
    input  input_45;
    input  input_46;
    input  input_47;
    input  input_48;
    input  input_49;
    input  input_50;
    input  input_51;
    input  input_52;
    input  input_53;
    input  input_54;
    input  input_55;
    input [5:0] sel;
    reg  result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      default : begin
        result = input_55;
      end
    endcase
    MUX_s_1_56_2 = result;
  end
  endfunction


  function automatic [1023:0] MUX_v_1024_2_2;
    input [1023:0] input_0;
    input [1023:0] input_1;
    input  sel;
    reg [1023:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_1024_2_2 = result;
  end
  endfunction


  function automatic [13:0] MUX_v_14_2_2;
    input [13:0] input_0;
    input [13:0] input_1;
    input  sel;
    reg [13:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_14_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_64_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [15:0] input_25;
    input [15:0] input_26;
    input [15:0] input_27;
    input [15:0] input_28;
    input [15:0] input_29;
    input [15:0] input_30;
    input [15:0] input_31;
    input [15:0] input_32;
    input [15:0] input_33;
    input [15:0] input_34;
    input [15:0] input_35;
    input [15:0] input_36;
    input [15:0] input_37;
    input [15:0] input_38;
    input [15:0] input_39;
    input [15:0] input_40;
    input [15:0] input_41;
    input [15:0] input_42;
    input [15:0] input_43;
    input [15:0] input_44;
    input [15:0] input_45;
    input [15:0] input_46;
    input [15:0] input_47;
    input [15:0] input_48;
    input [15:0] input_49;
    input [15:0] input_50;
    input [15:0] input_51;
    input [15:0] input_52;
    input [15:0] input_53;
    input [15:0] input_54;
    input [15:0] input_55;
    input [15:0] input_56;
    input [15:0] input_57;
    input [15:0] input_58;
    input [15:0] input_59;
    input [15:0] input_60;
    input [15:0] input_61;
    input [15:0] input_62;
    input [15:0] input_63;
    input [5:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      6'b000000 : begin
        result = input_0;
      end
      6'b000001 : begin
        result = input_1;
      end
      6'b000010 : begin
        result = input_2;
      end
      6'b000011 : begin
        result = input_3;
      end
      6'b000100 : begin
        result = input_4;
      end
      6'b000101 : begin
        result = input_5;
      end
      6'b000110 : begin
        result = input_6;
      end
      6'b000111 : begin
        result = input_7;
      end
      6'b001000 : begin
        result = input_8;
      end
      6'b001001 : begin
        result = input_9;
      end
      6'b001010 : begin
        result = input_10;
      end
      6'b001011 : begin
        result = input_11;
      end
      6'b001100 : begin
        result = input_12;
      end
      6'b001101 : begin
        result = input_13;
      end
      6'b001110 : begin
        result = input_14;
      end
      6'b001111 : begin
        result = input_15;
      end
      6'b010000 : begin
        result = input_16;
      end
      6'b010001 : begin
        result = input_17;
      end
      6'b010010 : begin
        result = input_18;
      end
      6'b010011 : begin
        result = input_19;
      end
      6'b010100 : begin
        result = input_20;
      end
      6'b010101 : begin
        result = input_21;
      end
      6'b010110 : begin
        result = input_22;
      end
      6'b010111 : begin
        result = input_23;
      end
      6'b011000 : begin
        result = input_24;
      end
      6'b011001 : begin
        result = input_25;
      end
      6'b011010 : begin
        result = input_26;
      end
      6'b011011 : begin
        result = input_27;
      end
      6'b011100 : begin
        result = input_28;
      end
      6'b011101 : begin
        result = input_29;
      end
      6'b011110 : begin
        result = input_30;
      end
      6'b011111 : begin
        result = input_31;
      end
      6'b100000 : begin
        result = input_32;
      end
      6'b100001 : begin
        result = input_33;
      end
      6'b100010 : begin
        result = input_34;
      end
      6'b100011 : begin
        result = input_35;
      end
      6'b100100 : begin
        result = input_36;
      end
      6'b100101 : begin
        result = input_37;
      end
      6'b100110 : begin
        result = input_38;
      end
      6'b100111 : begin
        result = input_39;
      end
      6'b101000 : begin
        result = input_40;
      end
      6'b101001 : begin
        result = input_41;
      end
      6'b101010 : begin
        result = input_42;
      end
      6'b101011 : begin
        result = input_43;
      end
      6'b101100 : begin
        result = input_44;
      end
      6'b101101 : begin
        result = input_45;
      end
      6'b101110 : begin
        result = input_46;
      end
      6'b101111 : begin
        result = input_47;
      end
      6'b110000 : begin
        result = input_48;
      end
      6'b110001 : begin
        result = input_49;
      end
      6'b110010 : begin
        result = input_50;
      end
      6'b110011 : begin
        result = input_51;
      end
      6'b110100 : begin
        result = input_52;
      end
      6'b110101 : begin
        result = input_53;
      end
      6'b110110 : begin
        result = input_54;
      end
      6'b110111 : begin
        result = input_55;
      end
      6'b111000 : begin
        result = input_56;
      end
      6'b111001 : begin
        result = input_57;
      end
      6'b111010 : begin
        result = input_58;
      end
      6'b111011 : begin
        result = input_59;
      end
      6'b111100 : begin
        result = input_60;
      end
      6'b111101 : begin
        result = input_61;
      end
      6'b111110 : begin
        result = input_62;
      end
      default : begin
        result = input_63;
      end
    endcase
    MUX_v_16_64_2 = result;
  end
  endfunction


  function automatic [19:0] MUX_v_20_2_2;
    input [19:0] input_0;
    input [19:0] input_1;
    input  sel;
    reg [19:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_20_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_15_1_14;
    input [14:0] vector;
    reg [14:0] tmp;
  begin
    tmp = vector >> 14;
    readslicef_15_1_14 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_22_1_21;
    input [21:0] vector;
    reg [21:0] tmp;
  begin
    tmp = vector >> 21;
    readslicef_22_1_21 = tmp[0:0];
  end
  endfunction


  function automatic [13:0] conv_s2s_8_14 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_14 = {{6{vector[7]}}, vector};
  end
  endfunction


  function automatic [14:0] conv_s2u_14_15 ;
    input [13:0]  vector ;
  begin
    conv_s2u_14_15 = {vector[13], vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_18_20 ;
    input [17:0]  vector ;
  begin
    conv_s2u_18_20 = {{2{vector[17]}}, vector};
  end
  endfunction


  function automatic [19:0] conv_s2u_19_20 ;
    input [18:0]  vector ;
  begin
    conv_s2u_19_20 = {vector[18], vector};
  end
  endfunction


  function automatic [20:0] conv_s2u_20_21 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_21 = {vector[19], vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_20_22 ;
    input [19:0]  vector ;
  begin
    conv_s2u_20_22 = {{2{vector[19]}}, vector};
  end
  endfunction


  function automatic [21:0] conv_s2u_21_22 ;
    input [20:0]  vector ;
  begin
    conv_s2u_21_22 = {vector[20], vector};
  end
  endfunction


  function automatic [3:0] conv_u2s_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2s_6_7 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Filter
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Filter (
  clk, rst, arst_n, head, length, dim, q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy,
      k_chan1_rsc_dat, k_chan1_rsc_vld, k_chan1_rsc_rdy, v_chan1_rsc_dat, v_chan1_rsc_vld,
      v_chan1_rsc_rdy, q_chan2_rsc_dat, q_chan2_rsc_vld, q_chan2_rsc_rdy, k_chan2_rsc_dat,
      k_chan2_rsc_vld, k_chan2_rsc_rdy, v_chan2_rsc_dat, v_chan2_rsc_vld, v_chan2_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [1023:0] q_chan1_rsc_dat;
  input q_chan1_rsc_vld;
  output q_chan1_rsc_rdy;
  input [1023:0] k_chan1_rsc_dat;
  input k_chan1_rsc_vld;
  output k_chan1_rsc_rdy;
  input [1023:0] v_chan1_rsc_dat;
  input v_chan1_rsc_vld;
  output v_chan1_rsc_rdy;
  output [1023:0] q_chan2_rsc_dat;
  output q_chan2_rsc_vld;
  input q_chan2_rsc_rdy;
  output [1023:0] k_chan2_rsc_dat;
  output k_chan2_rsc_vld;
  input k_chan2_rsc_rdy;
  output [1023:0] v_chan2_rsc_dat;
  output v_chan2_rsc_vld;
  input v_chan2_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ATTENTION_IP_Attention_Filter_run ATTENTION_IP_Attention_Filter_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .q_chan1_rsc_dat(q_chan1_rsc_dat),
      .q_chan1_rsc_vld(q_chan1_rsc_vld),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy),
      .k_chan1_rsc_dat(k_chan1_rsc_dat),
      .k_chan1_rsc_vld(k_chan1_rsc_vld),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy),
      .v_chan1_rsc_dat(v_chan1_rsc_dat),
      .v_chan1_rsc_vld(v_chan1_rsc_vld),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy),
      .q_chan2_rsc_dat(q_chan2_rsc_dat),
      .q_chan2_rsc_vld(q_chan2_rsc_vld),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy),
      .k_chan2_rsc_dat(k_chan2_rsc_dat),
      .k_chan2_rsc_vld(k_chan2_rsc_vld),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy),
      .v_chan2_rsc_dat(v_chan2_rsc_dat),
      .v_chan2_rsc_vld(v_chan2_rsc_vld),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy)
    );
endmodule




//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_in_wait_coupled_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_coupled_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/ccs_ram_sync_1R1W.v 
module ccs_ram_sync_1R1W
#(
parameter data_width = 8,
parameter addr_width = 7,
parameter depth = 128
)(
	radr, wadr, d, we, re, clk, q
);

	input [addr_width-1:0] radr;
	input [addr_width-1:0] wadr;
	input [data_width-1:0] d;
	input we;
	input re;
	input clk;
	output[data_width-1:0] q;

   // synopsys translate_off
	reg [data_width-1:0] q;

	reg [data_width-1:0] mem [depth-1:0];
		
	always @(posedge clk) begin
		if (we) begin
			mem[wadr] <= d; // Write port
		end
		if (re) begin
			q <= mem[radr] ; // read port
		end
	end
   // synopsys translate_on

endmodule

//------> ../ATTENTION_IP_Attention_Buffer.v2/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   b08092@cad29.ee.ntu.edu.tw
//  Generated date: Wed Jun 12 20:08:23 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_8_16_14_10752_10752_16_5_gen
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_8_16_14_10752_10752_16_5_gen
    (
  we, d, wadr, q, re, radr, radr_d, wadr_d, d_d, we_d, re_d, q_d, port_0_r_ram_ir_internal_RMASK_B_d,
      port_1_w_ram_ir_internal_WMASK_B_d
);
  output we;
  output [15:0] d;
  output [13:0] wadr;
  input [15:0] q;
  output re;
  output [13:0] radr;
  input [13:0] radr_d;
  input [13:0] wadr_d;
  input [15:0] d_d;
  input we_d;
  input re_d;
  output [15:0] q_d;
  input port_0_r_ram_ir_internal_RMASK_B_d;
  input port_1_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign we = (port_1_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
  assign q_d = q;
  assign re = (port_0_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, LOOPK1_C_0_tr0, LOOPJ1_C_64_tr0, LOOPK2_C_65_tr0,
      LOOPK3_C_65_tr0, LOOPJ2_C_66_tr0, LOOPI1_C_0_tr0
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;
  input LOOPK1_C_0_tr0;
  input LOOPJ1_C_64_tr0;
  input LOOPK2_C_65_tr0;
  input LOOPK3_C_65_tr0;
  input LOOPJ2_C_66_tr0;
  input LOOPI1_C_0_tr0;


  // FSM State Type Declaration for ATTENTION_IP_Attention_Buffer_run_run_fsm_1
  parameter
    main_C_0 = 9'd0,
    LOOPK1_C_0 = 9'd1,
    LOOPJ1_C_0 = 9'd2,
    LOOPJ1_C_1 = 9'd3,
    LOOPJ1_C_2 = 9'd4,
    LOOPJ1_C_3 = 9'd5,
    LOOPJ1_C_4 = 9'd6,
    LOOPJ1_C_5 = 9'd7,
    LOOPJ1_C_6 = 9'd8,
    LOOPJ1_C_7 = 9'd9,
    LOOPJ1_C_8 = 9'd10,
    LOOPJ1_C_9 = 9'd11,
    LOOPJ1_C_10 = 9'd12,
    LOOPJ1_C_11 = 9'd13,
    LOOPJ1_C_12 = 9'd14,
    LOOPJ1_C_13 = 9'd15,
    LOOPJ1_C_14 = 9'd16,
    LOOPJ1_C_15 = 9'd17,
    LOOPJ1_C_16 = 9'd18,
    LOOPJ1_C_17 = 9'd19,
    LOOPJ1_C_18 = 9'd20,
    LOOPJ1_C_19 = 9'd21,
    LOOPJ1_C_20 = 9'd22,
    LOOPJ1_C_21 = 9'd23,
    LOOPJ1_C_22 = 9'd24,
    LOOPJ1_C_23 = 9'd25,
    LOOPJ1_C_24 = 9'd26,
    LOOPJ1_C_25 = 9'd27,
    LOOPJ1_C_26 = 9'd28,
    LOOPJ1_C_27 = 9'd29,
    LOOPJ1_C_28 = 9'd30,
    LOOPJ1_C_29 = 9'd31,
    LOOPJ1_C_30 = 9'd32,
    LOOPJ1_C_31 = 9'd33,
    LOOPJ1_C_32 = 9'd34,
    LOOPJ1_C_33 = 9'd35,
    LOOPJ1_C_34 = 9'd36,
    LOOPJ1_C_35 = 9'd37,
    LOOPJ1_C_36 = 9'd38,
    LOOPJ1_C_37 = 9'd39,
    LOOPJ1_C_38 = 9'd40,
    LOOPJ1_C_39 = 9'd41,
    LOOPJ1_C_40 = 9'd42,
    LOOPJ1_C_41 = 9'd43,
    LOOPJ1_C_42 = 9'd44,
    LOOPJ1_C_43 = 9'd45,
    LOOPJ1_C_44 = 9'd46,
    LOOPJ1_C_45 = 9'd47,
    LOOPJ1_C_46 = 9'd48,
    LOOPJ1_C_47 = 9'd49,
    LOOPJ1_C_48 = 9'd50,
    LOOPJ1_C_49 = 9'd51,
    LOOPJ1_C_50 = 9'd52,
    LOOPJ1_C_51 = 9'd53,
    LOOPJ1_C_52 = 9'd54,
    LOOPJ1_C_53 = 9'd55,
    LOOPJ1_C_54 = 9'd56,
    LOOPJ1_C_55 = 9'd57,
    LOOPJ1_C_56 = 9'd58,
    LOOPJ1_C_57 = 9'd59,
    LOOPJ1_C_58 = 9'd60,
    LOOPJ1_C_59 = 9'd61,
    LOOPJ1_C_60 = 9'd62,
    LOOPJ1_C_61 = 9'd63,
    LOOPJ1_C_62 = 9'd64,
    LOOPJ1_C_63 = 9'd65,
    LOOPJ1_C_64 = 9'd66,
    LOOPJ2_C_0 = 9'd67,
    LOOPJ2_C_1 = 9'd68,
    LOOPJ2_C_2 = 9'd69,
    LOOPJ2_C_3 = 9'd70,
    LOOPJ2_C_4 = 9'd71,
    LOOPJ2_C_5 = 9'd72,
    LOOPJ2_C_6 = 9'd73,
    LOOPJ2_C_7 = 9'd74,
    LOOPJ2_C_8 = 9'd75,
    LOOPJ2_C_9 = 9'd76,
    LOOPJ2_C_10 = 9'd77,
    LOOPJ2_C_11 = 9'd78,
    LOOPJ2_C_12 = 9'd79,
    LOOPJ2_C_13 = 9'd80,
    LOOPJ2_C_14 = 9'd81,
    LOOPJ2_C_15 = 9'd82,
    LOOPJ2_C_16 = 9'd83,
    LOOPJ2_C_17 = 9'd84,
    LOOPJ2_C_18 = 9'd85,
    LOOPJ2_C_19 = 9'd86,
    LOOPJ2_C_20 = 9'd87,
    LOOPJ2_C_21 = 9'd88,
    LOOPJ2_C_22 = 9'd89,
    LOOPJ2_C_23 = 9'd90,
    LOOPJ2_C_24 = 9'd91,
    LOOPJ2_C_25 = 9'd92,
    LOOPJ2_C_26 = 9'd93,
    LOOPJ2_C_27 = 9'd94,
    LOOPJ2_C_28 = 9'd95,
    LOOPJ2_C_29 = 9'd96,
    LOOPJ2_C_30 = 9'd97,
    LOOPJ2_C_31 = 9'd98,
    LOOPJ2_C_32 = 9'd99,
    LOOPJ2_C_33 = 9'd100,
    LOOPJ2_C_34 = 9'd101,
    LOOPJ2_C_35 = 9'd102,
    LOOPJ2_C_36 = 9'd103,
    LOOPJ2_C_37 = 9'd104,
    LOOPJ2_C_38 = 9'd105,
    LOOPJ2_C_39 = 9'd106,
    LOOPJ2_C_40 = 9'd107,
    LOOPJ2_C_41 = 9'd108,
    LOOPJ2_C_42 = 9'd109,
    LOOPJ2_C_43 = 9'd110,
    LOOPJ2_C_44 = 9'd111,
    LOOPJ2_C_45 = 9'd112,
    LOOPJ2_C_46 = 9'd113,
    LOOPJ2_C_47 = 9'd114,
    LOOPJ2_C_48 = 9'd115,
    LOOPJ2_C_49 = 9'd116,
    LOOPJ2_C_50 = 9'd117,
    LOOPJ2_C_51 = 9'd118,
    LOOPJ2_C_52 = 9'd119,
    LOOPJ2_C_53 = 9'd120,
    LOOPJ2_C_54 = 9'd121,
    LOOPJ2_C_55 = 9'd122,
    LOOPJ2_C_56 = 9'd123,
    LOOPJ2_C_57 = 9'd124,
    LOOPJ2_C_58 = 9'd125,
    LOOPJ2_C_59 = 9'd126,
    LOOPJ2_C_60 = 9'd127,
    LOOPJ2_C_61 = 9'd128,
    LOOPJ2_C_62 = 9'd129,
    LOOPJ2_C_63 = 9'd130,
    LOOPJ2_C_64 = 9'd131,
    LOOPJ2_C_65 = 9'd132,
    LOOPK2_C_0 = 9'd133,
    LOOPK2_C_1 = 9'd134,
    LOOPK2_C_2 = 9'd135,
    LOOPK2_C_3 = 9'd136,
    LOOPK2_C_4 = 9'd137,
    LOOPK2_C_5 = 9'd138,
    LOOPK2_C_6 = 9'd139,
    LOOPK2_C_7 = 9'd140,
    LOOPK2_C_8 = 9'd141,
    LOOPK2_C_9 = 9'd142,
    LOOPK2_C_10 = 9'd143,
    LOOPK2_C_11 = 9'd144,
    LOOPK2_C_12 = 9'd145,
    LOOPK2_C_13 = 9'd146,
    LOOPK2_C_14 = 9'd147,
    LOOPK2_C_15 = 9'd148,
    LOOPK2_C_16 = 9'd149,
    LOOPK2_C_17 = 9'd150,
    LOOPK2_C_18 = 9'd151,
    LOOPK2_C_19 = 9'd152,
    LOOPK2_C_20 = 9'd153,
    LOOPK2_C_21 = 9'd154,
    LOOPK2_C_22 = 9'd155,
    LOOPK2_C_23 = 9'd156,
    LOOPK2_C_24 = 9'd157,
    LOOPK2_C_25 = 9'd158,
    LOOPK2_C_26 = 9'd159,
    LOOPK2_C_27 = 9'd160,
    LOOPK2_C_28 = 9'd161,
    LOOPK2_C_29 = 9'd162,
    LOOPK2_C_30 = 9'd163,
    LOOPK2_C_31 = 9'd164,
    LOOPK2_C_32 = 9'd165,
    LOOPK2_C_33 = 9'd166,
    LOOPK2_C_34 = 9'd167,
    LOOPK2_C_35 = 9'd168,
    LOOPK2_C_36 = 9'd169,
    LOOPK2_C_37 = 9'd170,
    LOOPK2_C_38 = 9'd171,
    LOOPK2_C_39 = 9'd172,
    LOOPK2_C_40 = 9'd173,
    LOOPK2_C_41 = 9'd174,
    LOOPK2_C_42 = 9'd175,
    LOOPK2_C_43 = 9'd176,
    LOOPK2_C_44 = 9'd177,
    LOOPK2_C_45 = 9'd178,
    LOOPK2_C_46 = 9'd179,
    LOOPK2_C_47 = 9'd180,
    LOOPK2_C_48 = 9'd181,
    LOOPK2_C_49 = 9'd182,
    LOOPK2_C_50 = 9'd183,
    LOOPK2_C_51 = 9'd184,
    LOOPK2_C_52 = 9'd185,
    LOOPK2_C_53 = 9'd186,
    LOOPK2_C_54 = 9'd187,
    LOOPK2_C_55 = 9'd188,
    LOOPK2_C_56 = 9'd189,
    LOOPK2_C_57 = 9'd190,
    LOOPK2_C_58 = 9'd191,
    LOOPK2_C_59 = 9'd192,
    LOOPK2_C_60 = 9'd193,
    LOOPK2_C_61 = 9'd194,
    LOOPK2_C_62 = 9'd195,
    LOOPK2_C_63 = 9'd196,
    LOOPK2_C_64 = 9'd197,
    LOOPK2_C_65 = 9'd198,
    LOOPK3_C_0 = 9'd199,
    LOOPK3_C_1 = 9'd200,
    LOOPK3_C_2 = 9'd201,
    LOOPK3_C_3 = 9'd202,
    LOOPK3_C_4 = 9'd203,
    LOOPK3_C_5 = 9'd204,
    LOOPK3_C_6 = 9'd205,
    LOOPK3_C_7 = 9'd206,
    LOOPK3_C_8 = 9'd207,
    LOOPK3_C_9 = 9'd208,
    LOOPK3_C_10 = 9'd209,
    LOOPK3_C_11 = 9'd210,
    LOOPK3_C_12 = 9'd211,
    LOOPK3_C_13 = 9'd212,
    LOOPK3_C_14 = 9'd213,
    LOOPK3_C_15 = 9'd214,
    LOOPK3_C_16 = 9'd215,
    LOOPK3_C_17 = 9'd216,
    LOOPK3_C_18 = 9'd217,
    LOOPK3_C_19 = 9'd218,
    LOOPK3_C_20 = 9'd219,
    LOOPK3_C_21 = 9'd220,
    LOOPK3_C_22 = 9'd221,
    LOOPK3_C_23 = 9'd222,
    LOOPK3_C_24 = 9'd223,
    LOOPK3_C_25 = 9'd224,
    LOOPK3_C_26 = 9'd225,
    LOOPK3_C_27 = 9'd226,
    LOOPK3_C_28 = 9'd227,
    LOOPK3_C_29 = 9'd228,
    LOOPK3_C_30 = 9'd229,
    LOOPK3_C_31 = 9'd230,
    LOOPK3_C_32 = 9'd231,
    LOOPK3_C_33 = 9'd232,
    LOOPK3_C_34 = 9'd233,
    LOOPK3_C_35 = 9'd234,
    LOOPK3_C_36 = 9'd235,
    LOOPK3_C_37 = 9'd236,
    LOOPK3_C_38 = 9'd237,
    LOOPK3_C_39 = 9'd238,
    LOOPK3_C_40 = 9'd239,
    LOOPK3_C_41 = 9'd240,
    LOOPK3_C_42 = 9'd241,
    LOOPK3_C_43 = 9'd242,
    LOOPK3_C_44 = 9'd243,
    LOOPK3_C_45 = 9'd244,
    LOOPK3_C_46 = 9'd245,
    LOOPK3_C_47 = 9'd246,
    LOOPK3_C_48 = 9'd247,
    LOOPK3_C_49 = 9'd248,
    LOOPK3_C_50 = 9'd249,
    LOOPK3_C_51 = 9'd250,
    LOOPK3_C_52 = 9'd251,
    LOOPK3_C_53 = 9'd252,
    LOOPK3_C_54 = 9'd253,
    LOOPK3_C_55 = 9'd254,
    LOOPK3_C_56 = 9'd255,
    LOOPK3_C_57 = 9'd256,
    LOOPK3_C_58 = 9'd257,
    LOOPK3_C_59 = 9'd258,
    LOOPK3_C_60 = 9'd259,
    LOOPK3_C_61 = 9'd260,
    LOOPK3_C_62 = 9'd261,
    LOOPK3_C_63 = 9'd262,
    LOOPK3_C_64 = 9'd263,
    LOOPK3_C_65 = 9'd264,
    LOOPJ2_C_66 = 9'd265,
    LOOPI1_C_0 = 9'd266,
    main_C_1 = 9'd267;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ATTENTION_IP_Attention_Buffer_run_run_fsm_1
    case (state_var)
      LOOPK1_C_0 : begin
        fsm_output = 9'b000000001;
        if ( LOOPK1_C_0_tr0 ) begin
          state_var_NS = LOOPJ1_C_0;
        end
        else begin
          state_var_NS = LOOPK1_C_0;
        end
      end
      LOOPJ1_C_0 : begin
        fsm_output = 9'b000000010;
        state_var_NS = LOOPJ1_C_1;
      end
      LOOPJ1_C_1 : begin
        fsm_output = 9'b000000011;
        state_var_NS = LOOPJ1_C_2;
      end
      LOOPJ1_C_2 : begin
        fsm_output = 9'b000000100;
        state_var_NS = LOOPJ1_C_3;
      end
      LOOPJ1_C_3 : begin
        fsm_output = 9'b000000101;
        state_var_NS = LOOPJ1_C_4;
      end
      LOOPJ1_C_4 : begin
        fsm_output = 9'b000000110;
        state_var_NS = LOOPJ1_C_5;
      end
      LOOPJ1_C_5 : begin
        fsm_output = 9'b000000111;
        state_var_NS = LOOPJ1_C_6;
      end
      LOOPJ1_C_6 : begin
        fsm_output = 9'b000001000;
        state_var_NS = LOOPJ1_C_7;
      end
      LOOPJ1_C_7 : begin
        fsm_output = 9'b000001001;
        state_var_NS = LOOPJ1_C_8;
      end
      LOOPJ1_C_8 : begin
        fsm_output = 9'b000001010;
        state_var_NS = LOOPJ1_C_9;
      end
      LOOPJ1_C_9 : begin
        fsm_output = 9'b000001011;
        state_var_NS = LOOPJ1_C_10;
      end
      LOOPJ1_C_10 : begin
        fsm_output = 9'b000001100;
        state_var_NS = LOOPJ1_C_11;
      end
      LOOPJ1_C_11 : begin
        fsm_output = 9'b000001101;
        state_var_NS = LOOPJ1_C_12;
      end
      LOOPJ1_C_12 : begin
        fsm_output = 9'b000001110;
        state_var_NS = LOOPJ1_C_13;
      end
      LOOPJ1_C_13 : begin
        fsm_output = 9'b000001111;
        state_var_NS = LOOPJ1_C_14;
      end
      LOOPJ1_C_14 : begin
        fsm_output = 9'b000010000;
        state_var_NS = LOOPJ1_C_15;
      end
      LOOPJ1_C_15 : begin
        fsm_output = 9'b000010001;
        state_var_NS = LOOPJ1_C_16;
      end
      LOOPJ1_C_16 : begin
        fsm_output = 9'b000010010;
        state_var_NS = LOOPJ1_C_17;
      end
      LOOPJ1_C_17 : begin
        fsm_output = 9'b000010011;
        state_var_NS = LOOPJ1_C_18;
      end
      LOOPJ1_C_18 : begin
        fsm_output = 9'b000010100;
        state_var_NS = LOOPJ1_C_19;
      end
      LOOPJ1_C_19 : begin
        fsm_output = 9'b000010101;
        state_var_NS = LOOPJ1_C_20;
      end
      LOOPJ1_C_20 : begin
        fsm_output = 9'b000010110;
        state_var_NS = LOOPJ1_C_21;
      end
      LOOPJ1_C_21 : begin
        fsm_output = 9'b000010111;
        state_var_NS = LOOPJ1_C_22;
      end
      LOOPJ1_C_22 : begin
        fsm_output = 9'b000011000;
        state_var_NS = LOOPJ1_C_23;
      end
      LOOPJ1_C_23 : begin
        fsm_output = 9'b000011001;
        state_var_NS = LOOPJ1_C_24;
      end
      LOOPJ1_C_24 : begin
        fsm_output = 9'b000011010;
        state_var_NS = LOOPJ1_C_25;
      end
      LOOPJ1_C_25 : begin
        fsm_output = 9'b000011011;
        state_var_NS = LOOPJ1_C_26;
      end
      LOOPJ1_C_26 : begin
        fsm_output = 9'b000011100;
        state_var_NS = LOOPJ1_C_27;
      end
      LOOPJ1_C_27 : begin
        fsm_output = 9'b000011101;
        state_var_NS = LOOPJ1_C_28;
      end
      LOOPJ1_C_28 : begin
        fsm_output = 9'b000011110;
        state_var_NS = LOOPJ1_C_29;
      end
      LOOPJ1_C_29 : begin
        fsm_output = 9'b000011111;
        state_var_NS = LOOPJ1_C_30;
      end
      LOOPJ1_C_30 : begin
        fsm_output = 9'b000100000;
        state_var_NS = LOOPJ1_C_31;
      end
      LOOPJ1_C_31 : begin
        fsm_output = 9'b000100001;
        state_var_NS = LOOPJ1_C_32;
      end
      LOOPJ1_C_32 : begin
        fsm_output = 9'b000100010;
        state_var_NS = LOOPJ1_C_33;
      end
      LOOPJ1_C_33 : begin
        fsm_output = 9'b000100011;
        state_var_NS = LOOPJ1_C_34;
      end
      LOOPJ1_C_34 : begin
        fsm_output = 9'b000100100;
        state_var_NS = LOOPJ1_C_35;
      end
      LOOPJ1_C_35 : begin
        fsm_output = 9'b000100101;
        state_var_NS = LOOPJ1_C_36;
      end
      LOOPJ1_C_36 : begin
        fsm_output = 9'b000100110;
        state_var_NS = LOOPJ1_C_37;
      end
      LOOPJ1_C_37 : begin
        fsm_output = 9'b000100111;
        state_var_NS = LOOPJ1_C_38;
      end
      LOOPJ1_C_38 : begin
        fsm_output = 9'b000101000;
        state_var_NS = LOOPJ1_C_39;
      end
      LOOPJ1_C_39 : begin
        fsm_output = 9'b000101001;
        state_var_NS = LOOPJ1_C_40;
      end
      LOOPJ1_C_40 : begin
        fsm_output = 9'b000101010;
        state_var_NS = LOOPJ1_C_41;
      end
      LOOPJ1_C_41 : begin
        fsm_output = 9'b000101011;
        state_var_NS = LOOPJ1_C_42;
      end
      LOOPJ1_C_42 : begin
        fsm_output = 9'b000101100;
        state_var_NS = LOOPJ1_C_43;
      end
      LOOPJ1_C_43 : begin
        fsm_output = 9'b000101101;
        state_var_NS = LOOPJ1_C_44;
      end
      LOOPJ1_C_44 : begin
        fsm_output = 9'b000101110;
        state_var_NS = LOOPJ1_C_45;
      end
      LOOPJ1_C_45 : begin
        fsm_output = 9'b000101111;
        state_var_NS = LOOPJ1_C_46;
      end
      LOOPJ1_C_46 : begin
        fsm_output = 9'b000110000;
        state_var_NS = LOOPJ1_C_47;
      end
      LOOPJ1_C_47 : begin
        fsm_output = 9'b000110001;
        state_var_NS = LOOPJ1_C_48;
      end
      LOOPJ1_C_48 : begin
        fsm_output = 9'b000110010;
        state_var_NS = LOOPJ1_C_49;
      end
      LOOPJ1_C_49 : begin
        fsm_output = 9'b000110011;
        state_var_NS = LOOPJ1_C_50;
      end
      LOOPJ1_C_50 : begin
        fsm_output = 9'b000110100;
        state_var_NS = LOOPJ1_C_51;
      end
      LOOPJ1_C_51 : begin
        fsm_output = 9'b000110101;
        state_var_NS = LOOPJ1_C_52;
      end
      LOOPJ1_C_52 : begin
        fsm_output = 9'b000110110;
        state_var_NS = LOOPJ1_C_53;
      end
      LOOPJ1_C_53 : begin
        fsm_output = 9'b000110111;
        state_var_NS = LOOPJ1_C_54;
      end
      LOOPJ1_C_54 : begin
        fsm_output = 9'b000111000;
        state_var_NS = LOOPJ1_C_55;
      end
      LOOPJ1_C_55 : begin
        fsm_output = 9'b000111001;
        state_var_NS = LOOPJ1_C_56;
      end
      LOOPJ1_C_56 : begin
        fsm_output = 9'b000111010;
        state_var_NS = LOOPJ1_C_57;
      end
      LOOPJ1_C_57 : begin
        fsm_output = 9'b000111011;
        state_var_NS = LOOPJ1_C_58;
      end
      LOOPJ1_C_58 : begin
        fsm_output = 9'b000111100;
        state_var_NS = LOOPJ1_C_59;
      end
      LOOPJ1_C_59 : begin
        fsm_output = 9'b000111101;
        state_var_NS = LOOPJ1_C_60;
      end
      LOOPJ1_C_60 : begin
        fsm_output = 9'b000111110;
        state_var_NS = LOOPJ1_C_61;
      end
      LOOPJ1_C_61 : begin
        fsm_output = 9'b000111111;
        state_var_NS = LOOPJ1_C_62;
      end
      LOOPJ1_C_62 : begin
        fsm_output = 9'b001000000;
        state_var_NS = LOOPJ1_C_63;
      end
      LOOPJ1_C_63 : begin
        fsm_output = 9'b001000001;
        state_var_NS = LOOPJ1_C_64;
      end
      LOOPJ1_C_64 : begin
        fsm_output = 9'b001000010;
        if ( LOOPJ1_C_64_tr0 ) begin
          state_var_NS = LOOPJ2_C_0;
        end
        else begin
          state_var_NS = LOOPK1_C_0;
        end
      end
      LOOPJ2_C_0 : begin
        fsm_output = 9'b001000011;
        state_var_NS = LOOPJ2_C_1;
      end
      LOOPJ2_C_1 : begin
        fsm_output = 9'b001000100;
        state_var_NS = LOOPJ2_C_2;
      end
      LOOPJ2_C_2 : begin
        fsm_output = 9'b001000101;
        state_var_NS = LOOPJ2_C_3;
      end
      LOOPJ2_C_3 : begin
        fsm_output = 9'b001000110;
        state_var_NS = LOOPJ2_C_4;
      end
      LOOPJ2_C_4 : begin
        fsm_output = 9'b001000111;
        state_var_NS = LOOPJ2_C_5;
      end
      LOOPJ2_C_5 : begin
        fsm_output = 9'b001001000;
        state_var_NS = LOOPJ2_C_6;
      end
      LOOPJ2_C_6 : begin
        fsm_output = 9'b001001001;
        state_var_NS = LOOPJ2_C_7;
      end
      LOOPJ2_C_7 : begin
        fsm_output = 9'b001001010;
        state_var_NS = LOOPJ2_C_8;
      end
      LOOPJ2_C_8 : begin
        fsm_output = 9'b001001011;
        state_var_NS = LOOPJ2_C_9;
      end
      LOOPJ2_C_9 : begin
        fsm_output = 9'b001001100;
        state_var_NS = LOOPJ2_C_10;
      end
      LOOPJ2_C_10 : begin
        fsm_output = 9'b001001101;
        state_var_NS = LOOPJ2_C_11;
      end
      LOOPJ2_C_11 : begin
        fsm_output = 9'b001001110;
        state_var_NS = LOOPJ2_C_12;
      end
      LOOPJ2_C_12 : begin
        fsm_output = 9'b001001111;
        state_var_NS = LOOPJ2_C_13;
      end
      LOOPJ2_C_13 : begin
        fsm_output = 9'b001010000;
        state_var_NS = LOOPJ2_C_14;
      end
      LOOPJ2_C_14 : begin
        fsm_output = 9'b001010001;
        state_var_NS = LOOPJ2_C_15;
      end
      LOOPJ2_C_15 : begin
        fsm_output = 9'b001010010;
        state_var_NS = LOOPJ2_C_16;
      end
      LOOPJ2_C_16 : begin
        fsm_output = 9'b001010011;
        state_var_NS = LOOPJ2_C_17;
      end
      LOOPJ2_C_17 : begin
        fsm_output = 9'b001010100;
        state_var_NS = LOOPJ2_C_18;
      end
      LOOPJ2_C_18 : begin
        fsm_output = 9'b001010101;
        state_var_NS = LOOPJ2_C_19;
      end
      LOOPJ2_C_19 : begin
        fsm_output = 9'b001010110;
        state_var_NS = LOOPJ2_C_20;
      end
      LOOPJ2_C_20 : begin
        fsm_output = 9'b001010111;
        state_var_NS = LOOPJ2_C_21;
      end
      LOOPJ2_C_21 : begin
        fsm_output = 9'b001011000;
        state_var_NS = LOOPJ2_C_22;
      end
      LOOPJ2_C_22 : begin
        fsm_output = 9'b001011001;
        state_var_NS = LOOPJ2_C_23;
      end
      LOOPJ2_C_23 : begin
        fsm_output = 9'b001011010;
        state_var_NS = LOOPJ2_C_24;
      end
      LOOPJ2_C_24 : begin
        fsm_output = 9'b001011011;
        state_var_NS = LOOPJ2_C_25;
      end
      LOOPJ2_C_25 : begin
        fsm_output = 9'b001011100;
        state_var_NS = LOOPJ2_C_26;
      end
      LOOPJ2_C_26 : begin
        fsm_output = 9'b001011101;
        state_var_NS = LOOPJ2_C_27;
      end
      LOOPJ2_C_27 : begin
        fsm_output = 9'b001011110;
        state_var_NS = LOOPJ2_C_28;
      end
      LOOPJ2_C_28 : begin
        fsm_output = 9'b001011111;
        state_var_NS = LOOPJ2_C_29;
      end
      LOOPJ2_C_29 : begin
        fsm_output = 9'b001100000;
        state_var_NS = LOOPJ2_C_30;
      end
      LOOPJ2_C_30 : begin
        fsm_output = 9'b001100001;
        state_var_NS = LOOPJ2_C_31;
      end
      LOOPJ2_C_31 : begin
        fsm_output = 9'b001100010;
        state_var_NS = LOOPJ2_C_32;
      end
      LOOPJ2_C_32 : begin
        fsm_output = 9'b001100011;
        state_var_NS = LOOPJ2_C_33;
      end
      LOOPJ2_C_33 : begin
        fsm_output = 9'b001100100;
        state_var_NS = LOOPJ2_C_34;
      end
      LOOPJ2_C_34 : begin
        fsm_output = 9'b001100101;
        state_var_NS = LOOPJ2_C_35;
      end
      LOOPJ2_C_35 : begin
        fsm_output = 9'b001100110;
        state_var_NS = LOOPJ2_C_36;
      end
      LOOPJ2_C_36 : begin
        fsm_output = 9'b001100111;
        state_var_NS = LOOPJ2_C_37;
      end
      LOOPJ2_C_37 : begin
        fsm_output = 9'b001101000;
        state_var_NS = LOOPJ2_C_38;
      end
      LOOPJ2_C_38 : begin
        fsm_output = 9'b001101001;
        state_var_NS = LOOPJ2_C_39;
      end
      LOOPJ2_C_39 : begin
        fsm_output = 9'b001101010;
        state_var_NS = LOOPJ2_C_40;
      end
      LOOPJ2_C_40 : begin
        fsm_output = 9'b001101011;
        state_var_NS = LOOPJ2_C_41;
      end
      LOOPJ2_C_41 : begin
        fsm_output = 9'b001101100;
        state_var_NS = LOOPJ2_C_42;
      end
      LOOPJ2_C_42 : begin
        fsm_output = 9'b001101101;
        state_var_NS = LOOPJ2_C_43;
      end
      LOOPJ2_C_43 : begin
        fsm_output = 9'b001101110;
        state_var_NS = LOOPJ2_C_44;
      end
      LOOPJ2_C_44 : begin
        fsm_output = 9'b001101111;
        state_var_NS = LOOPJ2_C_45;
      end
      LOOPJ2_C_45 : begin
        fsm_output = 9'b001110000;
        state_var_NS = LOOPJ2_C_46;
      end
      LOOPJ2_C_46 : begin
        fsm_output = 9'b001110001;
        state_var_NS = LOOPJ2_C_47;
      end
      LOOPJ2_C_47 : begin
        fsm_output = 9'b001110010;
        state_var_NS = LOOPJ2_C_48;
      end
      LOOPJ2_C_48 : begin
        fsm_output = 9'b001110011;
        state_var_NS = LOOPJ2_C_49;
      end
      LOOPJ2_C_49 : begin
        fsm_output = 9'b001110100;
        state_var_NS = LOOPJ2_C_50;
      end
      LOOPJ2_C_50 : begin
        fsm_output = 9'b001110101;
        state_var_NS = LOOPJ2_C_51;
      end
      LOOPJ2_C_51 : begin
        fsm_output = 9'b001110110;
        state_var_NS = LOOPJ2_C_52;
      end
      LOOPJ2_C_52 : begin
        fsm_output = 9'b001110111;
        state_var_NS = LOOPJ2_C_53;
      end
      LOOPJ2_C_53 : begin
        fsm_output = 9'b001111000;
        state_var_NS = LOOPJ2_C_54;
      end
      LOOPJ2_C_54 : begin
        fsm_output = 9'b001111001;
        state_var_NS = LOOPJ2_C_55;
      end
      LOOPJ2_C_55 : begin
        fsm_output = 9'b001111010;
        state_var_NS = LOOPJ2_C_56;
      end
      LOOPJ2_C_56 : begin
        fsm_output = 9'b001111011;
        state_var_NS = LOOPJ2_C_57;
      end
      LOOPJ2_C_57 : begin
        fsm_output = 9'b001111100;
        state_var_NS = LOOPJ2_C_58;
      end
      LOOPJ2_C_58 : begin
        fsm_output = 9'b001111101;
        state_var_NS = LOOPJ2_C_59;
      end
      LOOPJ2_C_59 : begin
        fsm_output = 9'b001111110;
        state_var_NS = LOOPJ2_C_60;
      end
      LOOPJ2_C_60 : begin
        fsm_output = 9'b001111111;
        state_var_NS = LOOPJ2_C_61;
      end
      LOOPJ2_C_61 : begin
        fsm_output = 9'b010000000;
        state_var_NS = LOOPJ2_C_62;
      end
      LOOPJ2_C_62 : begin
        fsm_output = 9'b010000001;
        state_var_NS = LOOPJ2_C_63;
      end
      LOOPJ2_C_63 : begin
        fsm_output = 9'b010000010;
        state_var_NS = LOOPJ2_C_64;
      end
      LOOPJ2_C_64 : begin
        fsm_output = 9'b010000011;
        state_var_NS = LOOPJ2_C_65;
      end
      LOOPJ2_C_65 : begin
        fsm_output = 9'b010000100;
        state_var_NS = LOOPK2_C_0;
      end
      LOOPK2_C_0 : begin
        fsm_output = 9'b010000101;
        state_var_NS = LOOPK2_C_1;
      end
      LOOPK2_C_1 : begin
        fsm_output = 9'b010000110;
        state_var_NS = LOOPK2_C_2;
      end
      LOOPK2_C_2 : begin
        fsm_output = 9'b010000111;
        state_var_NS = LOOPK2_C_3;
      end
      LOOPK2_C_3 : begin
        fsm_output = 9'b010001000;
        state_var_NS = LOOPK2_C_4;
      end
      LOOPK2_C_4 : begin
        fsm_output = 9'b010001001;
        state_var_NS = LOOPK2_C_5;
      end
      LOOPK2_C_5 : begin
        fsm_output = 9'b010001010;
        state_var_NS = LOOPK2_C_6;
      end
      LOOPK2_C_6 : begin
        fsm_output = 9'b010001011;
        state_var_NS = LOOPK2_C_7;
      end
      LOOPK2_C_7 : begin
        fsm_output = 9'b010001100;
        state_var_NS = LOOPK2_C_8;
      end
      LOOPK2_C_8 : begin
        fsm_output = 9'b010001101;
        state_var_NS = LOOPK2_C_9;
      end
      LOOPK2_C_9 : begin
        fsm_output = 9'b010001110;
        state_var_NS = LOOPK2_C_10;
      end
      LOOPK2_C_10 : begin
        fsm_output = 9'b010001111;
        state_var_NS = LOOPK2_C_11;
      end
      LOOPK2_C_11 : begin
        fsm_output = 9'b010010000;
        state_var_NS = LOOPK2_C_12;
      end
      LOOPK2_C_12 : begin
        fsm_output = 9'b010010001;
        state_var_NS = LOOPK2_C_13;
      end
      LOOPK2_C_13 : begin
        fsm_output = 9'b010010010;
        state_var_NS = LOOPK2_C_14;
      end
      LOOPK2_C_14 : begin
        fsm_output = 9'b010010011;
        state_var_NS = LOOPK2_C_15;
      end
      LOOPK2_C_15 : begin
        fsm_output = 9'b010010100;
        state_var_NS = LOOPK2_C_16;
      end
      LOOPK2_C_16 : begin
        fsm_output = 9'b010010101;
        state_var_NS = LOOPK2_C_17;
      end
      LOOPK2_C_17 : begin
        fsm_output = 9'b010010110;
        state_var_NS = LOOPK2_C_18;
      end
      LOOPK2_C_18 : begin
        fsm_output = 9'b010010111;
        state_var_NS = LOOPK2_C_19;
      end
      LOOPK2_C_19 : begin
        fsm_output = 9'b010011000;
        state_var_NS = LOOPK2_C_20;
      end
      LOOPK2_C_20 : begin
        fsm_output = 9'b010011001;
        state_var_NS = LOOPK2_C_21;
      end
      LOOPK2_C_21 : begin
        fsm_output = 9'b010011010;
        state_var_NS = LOOPK2_C_22;
      end
      LOOPK2_C_22 : begin
        fsm_output = 9'b010011011;
        state_var_NS = LOOPK2_C_23;
      end
      LOOPK2_C_23 : begin
        fsm_output = 9'b010011100;
        state_var_NS = LOOPK2_C_24;
      end
      LOOPK2_C_24 : begin
        fsm_output = 9'b010011101;
        state_var_NS = LOOPK2_C_25;
      end
      LOOPK2_C_25 : begin
        fsm_output = 9'b010011110;
        state_var_NS = LOOPK2_C_26;
      end
      LOOPK2_C_26 : begin
        fsm_output = 9'b010011111;
        state_var_NS = LOOPK2_C_27;
      end
      LOOPK2_C_27 : begin
        fsm_output = 9'b010100000;
        state_var_NS = LOOPK2_C_28;
      end
      LOOPK2_C_28 : begin
        fsm_output = 9'b010100001;
        state_var_NS = LOOPK2_C_29;
      end
      LOOPK2_C_29 : begin
        fsm_output = 9'b010100010;
        state_var_NS = LOOPK2_C_30;
      end
      LOOPK2_C_30 : begin
        fsm_output = 9'b010100011;
        state_var_NS = LOOPK2_C_31;
      end
      LOOPK2_C_31 : begin
        fsm_output = 9'b010100100;
        state_var_NS = LOOPK2_C_32;
      end
      LOOPK2_C_32 : begin
        fsm_output = 9'b010100101;
        state_var_NS = LOOPK2_C_33;
      end
      LOOPK2_C_33 : begin
        fsm_output = 9'b010100110;
        state_var_NS = LOOPK2_C_34;
      end
      LOOPK2_C_34 : begin
        fsm_output = 9'b010100111;
        state_var_NS = LOOPK2_C_35;
      end
      LOOPK2_C_35 : begin
        fsm_output = 9'b010101000;
        state_var_NS = LOOPK2_C_36;
      end
      LOOPK2_C_36 : begin
        fsm_output = 9'b010101001;
        state_var_NS = LOOPK2_C_37;
      end
      LOOPK2_C_37 : begin
        fsm_output = 9'b010101010;
        state_var_NS = LOOPK2_C_38;
      end
      LOOPK2_C_38 : begin
        fsm_output = 9'b010101011;
        state_var_NS = LOOPK2_C_39;
      end
      LOOPK2_C_39 : begin
        fsm_output = 9'b010101100;
        state_var_NS = LOOPK2_C_40;
      end
      LOOPK2_C_40 : begin
        fsm_output = 9'b010101101;
        state_var_NS = LOOPK2_C_41;
      end
      LOOPK2_C_41 : begin
        fsm_output = 9'b010101110;
        state_var_NS = LOOPK2_C_42;
      end
      LOOPK2_C_42 : begin
        fsm_output = 9'b010101111;
        state_var_NS = LOOPK2_C_43;
      end
      LOOPK2_C_43 : begin
        fsm_output = 9'b010110000;
        state_var_NS = LOOPK2_C_44;
      end
      LOOPK2_C_44 : begin
        fsm_output = 9'b010110001;
        state_var_NS = LOOPK2_C_45;
      end
      LOOPK2_C_45 : begin
        fsm_output = 9'b010110010;
        state_var_NS = LOOPK2_C_46;
      end
      LOOPK2_C_46 : begin
        fsm_output = 9'b010110011;
        state_var_NS = LOOPK2_C_47;
      end
      LOOPK2_C_47 : begin
        fsm_output = 9'b010110100;
        state_var_NS = LOOPK2_C_48;
      end
      LOOPK2_C_48 : begin
        fsm_output = 9'b010110101;
        state_var_NS = LOOPK2_C_49;
      end
      LOOPK2_C_49 : begin
        fsm_output = 9'b010110110;
        state_var_NS = LOOPK2_C_50;
      end
      LOOPK2_C_50 : begin
        fsm_output = 9'b010110111;
        state_var_NS = LOOPK2_C_51;
      end
      LOOPK2_C_51 : begin
        fsm_output = 9'b010111000;
        state_var_NS = LOOPK2_C_52;
      end
      LOOPK2_C_52 : begin
        fsm_output = 9'b010111001;
        state_var_NS = LOOPK2_C_53;
      end
      LOOPK2_C_53 : begin
        fsm_output = 9'b010111010;
        state_var_NS = LOOPK2_C_54;
      end
      LOOPK2_C_54 : begin
        fsm_output = 9'b010111011;
        state_var_NS = LOOPK2_C_55;
      end
      LOOPK2_C_55 : begin
        fsm_output = 9'b010111100;
        state_var_NS = LOOPK2_C_56;
      end
      LOOPK2_C_56 : begin
        fsm_output = 9'b010111101;
        state_var_NS = LOOPK2_C_57;
      end
      LOOPK2_C_57 : begin
        fsm_output = 9'b010111110;
        state_var_NS = LOOPK2_C_58;
      end
      LOOPK2_C_58 : begin
        fsm_output = 9'b010111111;
        state_var_NS = LOOPK2_C_59;
      end
      LOOPK2_C_59 : begin
        fsm_output = 9'b011000000;
        state_var_NS = LOOPK2_C_60;
      end
      LOOPK2_C_60 : begin
        fsm_output = 9'b011000001;
        state_var_NS = LOOPK2_C_61;
      end
      LOOPK2_C_61 : begin
        fsm_output = 9'b011000010;
        state_var_NS = LOOPK2_C_62;
      end
      LOOPK2_C_62 : begin
        fsm_output = 9'b011000011;
        state_var_NS = LOOPK2_C_63;
      end
      LOOPK2_C_63 : begin
        fsm_output = 9'b011000100;
        state_var_NS = LOOPK2_C_64;
      end
      LOOPK2_C_64 : begin
        fsm_output = 9'b011000101;
        state_var_NS = LOOPK2_C_65;
      end
      LOOPK2_C_65 : begin
        fsm_output = 9'b011000110;
        if ( LOOPK2_C_65_tr0 ) begin
          state_var_NS = LOOPK3_C_0;
        end
        else begin
          state_var_NS = LOOPK2_C_0;
        end
      end
      LOOPK3_C_0 : begin
        fsm_output = 9'b011000111;
        state_var_NS = LOOPK3_C_1;
      end
      LOOPK3_C_1 : begin
        fsm_output = 9'b011001000;
        state_var_NS = LOOPK3_C_2;
      end
      LOOPK3_C_2 : begin
        fsm_output = 9'b011001001;
        state_var_NS = LOOPK3_C_3;
      end
      LOOPK3_C_3 : begin
        fsm_output = 9'b011001010;
        state_var_NS = LOOPK3_C_4;
      end
      LOOPK3_C_4 : begin
        fsm_output = 9'b011001011;
        state_var_NS = LOOPK3_C_5;
      end
      LOOPK3_C_5 : begin
        fsm_output = 9'b011001100;
        state_var_NS = LOOPK3_C_6;
      end
      LOOPK3_C_6 : begin
        fsm_output = 9'b011001101;
        state_var_NS = LOOPK3_C_7;
      end
      LOOPK3_C_7 : begin
        fsm_output = 9'b011001110;
        state_var_NS = LOOPK3_C_8;
      end
      LOOPK3_C_8 : begin
        fsm_output = 9'b011001111;
        state_var_NS = LOOPK3_C_9;
      end
      LOOPK3_C_9 : begin
        fsm_output = 9'b011010000;
        state_var_NS = LOOPK3_C_10;
      end
      LOOPK3_C_10 : begin
        fsm_output = 9'b011010001;
        state_var_NS = LOOPK3_C_11;
      end
      LOOPK3_C_11 : begin
        fsm_output = 9'b011010010;
        state_var_NS = LOOPK3_C_12;
      end
      LOOPK3_C_12 : begin
        fsm_output = 9'b011010011;
        state_var_NS = LOOPK3_C_13;
      end
      LOOPK3_C_13 : begin
        fsm_output = 9'b011010100;
        state_var_NS = LOOPK3_C_14;
      end
      LOOPK3_C_14 : begin
        fsm_output = 9'b011010101;
        state_var_NS = LOOPK3_C_15;
      end
      LOOPK3_C_15 : begin
        fsm_output = 9'b011010110;
        state_var_NS = LOOPK3_C_16;
      end
      LOOPK3_C_16 : begin
        fsm_output = 9'b011010111;
        state_var_NS = LOOPK3_C_17;
      end
      LOOPK3_C_17 : begin
        fsm_output = 9'b011011000;
        state_var_NS = LOOPK3_C_18;
      end
      LOOPK3_C_18 : begin
        fsm_output = 9'b011011001;
        state_var_NS = LOOPK3_C_19;
      end
      LOOPK3_C_19 : begin
        fsm_output = 9'b011011010;
        state_var_NS = LOOPK3_C_20;
      end
      LOOPK3_C_20 : begin
        fsm_output = 9'b011011011;
        state_var_NS = LOOPK3_C_21;
      end
      LOOPK3_C_21 : begin
        fsm_output = 9'b011011100;
        state_var_NS = LOOPK3_C_22;
      end
      LOOPK3_C_22 : begin
        fsm_output = 9'b011011101;
        state_var_NS = LOOPK3_C_23;
      end
      LOOPK3_C_23 : begin
        fsm_output = 9'b011011110;
        state_var_NS = LOOPK3_C_24;
      end
      LOOPK3_C_24 : begin
        fsm_output = 9'b011011111;
        state_var_NS = LOOPK3_C_25;
      end
      LOOPK3_C_25 : begin
        fsm_output = 9'b011100000;
        state_var_NS = LOOPK3_C_26;
      end
      LOOPK3_C_26 : begin
        fsm_output = 9'b011100001;
        state_var_NS = LOOPK3_C_27;
      end
      LOOPK3_C_27 : begin
        fsm_output = 9'b011100010;
        state_var_NS = LOOPK3_C_28;
      end
      LOOPK3_C_28 : begin
        fsm_output = 9'b011100011;
        state_var_NS = LOOPK3_C_29;
      end
      LOOPK3_C_29 : begin
        fsm_output = 9'b011100100;
        state_var_NS = LOOPK3_C_30;
      end
      LOOPK3_C_30 : begin
        fsm_output = 9'b011100101;
        state_var_NS = LOOPK3_C_31;
      end
      LOOPK3_C_31 : begin
        fsm_output = 9'b011100110;
        state_var_NS = LOOPK3_C_32;
      end
      LOOPK3_C_32 : begin
        fsm_output = 9'b011100111;
        state_var_NS = LOOPK3_C_33;
      end
      LOOPK3_C_33 : begin
        fsm_output = 9'b011101000;
        state_var_NS = LOOPK3_C_34;
      end
      LOOPK3_C_34 : begin
        fsm_output = 9'b011101001;
        state_var_NS = LOOPK3_C_35;
      end
      LOOPK3_C_35 : begin
        fsm_output = 9'b011101010;
        state_var_NS = LOOPK3_C_36;
      end
      LOOPK3_C_36 : begin
        fsm_output = 9'b011101011;
        state_var_NS = LOOPK3_C_37;
      end
      LOOPK3_C_37 : begin
        fsm_output = 9'b011101100;
        state_var_NS = LOOPK3_C_38;
      end
      LOOPK3_C_38 : begin
        fsm_output = 9'b011101101;
        state_var_NS = LOOPK3_C_39;
      end
      LOOPK3_C_39 : begin
        fsm_output = 9'b011101110;
        state_var_NS = LOOPK3_C_40;
      end
      LOOPK3_C_40 : begin
        fsm_output = 9'b011101111;
        state_var_NS = LOOPK3_C_41;
      end
      LOOPK3_C_41 : begin
        fsm_output = 9'b011110000;
        state_var_NS = LOOPK3_C_42;
      end
      LOOPK3_C_42 : begin
        fsm_output = 9'b011110001;
        state_var_NS = LOOPK3_C_43;
      end
      LOOPK3_C_43 : begin
        fsm_output = 9'b011110010;
        state_var_NS = LOOPK3_C_44;
      end
      LOOPK3_C_44 : begin
        fsm_output = 9'b011110011;
        state_var_NS = LOOPK3_C_45;
      end
      LOOPK3_C_45 : begin
        fsm_output = 9'b011110100;
        state_var_NS = LOOPK3_C_46;
      end
      LOOPK3_C_46 : begin
        fsm_output = 9'b011110101;
        state_var_NS = LOOPK3_C_47;
      end
      LOOPK3_C_47 : begin
        fsm_output = 9'b011110110;
        state_var_NS = LOOPK3_C_48;
      end
      LOOPK3_C_48 : begin
        fsm_output = 9'b011110111;
        state_var_NS = LOOPK3_C_49;
      end
      LOOPK3_C_49 : begin
        fsm_output = 9'b011111000;
        state_var_NS = LOOPK3_C_50;
      end
      LOOPK3_C_50 : begin
        fsm_output = 9'b011111001;
        state_var_NS = LOOPK3_C_51;
      end
      LOOPK3_C_51 : begin
        fsm_output = 9'b011111010;
        state_var_NS = LOOPK3_C_52;
      end
      LOOPK3_C_52 : begin
        fsm_output = 9'b011111011;
        state_var_NS = LOOPK3_C_53;
      end
      LOOPK3_C_53 : begin
        fsm_output = 9'b011111100;
        state_var_NS = LOOPK3_C_54;
      end
      LOOPK3_C_54 : begin
        fsm_output = 9'b011111101;
        state_var_NS = LOOPK3_C_55;
      end
      LOOPK3_C_55 : begin
        fsm_output = 9'b011111110;
        state_var_NS = LOOPK3_C_56;
      end
      LOOPK3_C_56 : begin
        fsm_output = 9'b011111111;
        state_var_NS = LOOPK3_C_57;
      end
      LOOPK3_C_57 : begin
        fsm_output = 9'b100000000;
        state_var_NS = LOOPK3_C_58;
      end
      LOOPK3_C_58 : begin
        fsm_output = 9'b100000001;
        state_var_NS = LOOPK3_C_59;
      end
      LOOPK3_C_59 : begin
        fsm_output = 9'b100000010;
        state_var_NS = LOOPK3_C_60;
      end
      LOOPK3_C_60 : begin
        fsm_output = 9'b100000011;
        state_var_NS = LOOPK3_C_61;
      end
      LOOPK3_C_61 : begin
        fsm_output = 9'b100000100;
        state_var_NS = LOOPK3_C_62;
      end
      LOOPK3_C_62 : begin
        fsm_output = 9'b100000101;
        state_var_NS = LOOPK3_C_63;
      end
      LOOPK3_C_63 : begin
        fsm_output = 9'b100000110;
        state_var_NS = LOOPK3_C_64;
      end
      LOOPK3_C_64 : begin
        fsm_output = 9'b100000111;
        state_var_NS = LOOPK3_C_65;
      end
      LOOPK3_C_65 : begin
        fsm_output = 9'b100001000;
        if ( LOOPK3_C_65_tr0 ) begin
          state_var_NS = LOOPJ2_C_66;
        end
        else begin
          state_var_NS = LOOPK3_C_0;
        end
      end
      LOOPJ2_C_66 : begin
        fsm_output = 9'b100001001;
        if ( LOOPJ2_C_66_tr0 ) begin
          state_var_NS = LOOPI1_C_0;
        end
        else begin
          state_var_NS = LOOPJ2_C_0;
        end
      end
      LOOPI1_C_0 : begin
        fsm_output = 9'b100001010;
        if ( LOOPI1_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = LOOPK1_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 9'b100001011;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = LOOPK1_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_staller
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_staller (
  clk, rst, arst_n, run_wen, run_wten, din_chan_rsci_wen_comp, q_chan1_rsci_wen_comp,
      k_chan1_rsci_wen_comp, v_chan1_rsci_wen_comp
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  output run_wten;
  input din_chan_rsci_wen_comp;
  input q_chan1_rsci_wen_comp;
  input k_chan1_rsci_wen_comp;
  input v_chan1_rsci_wen_comp;


  // Interconnect Declarations
  reg run_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = din_chan_rsci_wen_comp & q_chan1_rsci_wen_comp & k_chan1_rsci_wen_comp
      & v_chan1_rsci_wen_comp;
  assign run_wten = run_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_wten_reg <= 1'b0;
    end
    else if ( rst ) begin
      run_wten_reg <= 1'b0;
    end
    else begin
      run_wten_reg <= ~ run_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_dp
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_dp
    (
  clk, rst, arst_n, pp_buf_data_rsci_q_d, pp_buf_data_rsci_q_d_mxwt, pp_buf_data_rsci_biwt_1,
      pp_buf_data_rsci_bdwt_2
);
  input clk;
  input rst;
  input arst_n;
  input [15:0] pp_buf_data_rsci_q_d;
  output [15:0] pp_buf_data_rsci_q_d_mxwt;
  input pp_buf_data_rsci_biwt_1;
  input pp_buf_data_rsci_bdwt_2;


  // Interconnect Declarations
  reg pp_buf_data_rsci_bcwt_1;
  reg [15:0] pp_buf_data_rsci_q_d_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign pp_buf_data_rsci_q_d_mxwt = MUX_v_16_2_2(pp_buf_data_rsci_q_d, pp_buf_data_rsci_q_d_bfwt,
      pp_buf_data_rsci_bcwt_1);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      pp_buf_data_rsci_bcwt_1 <= 1'b0;
    end
    else if ( rst ) begin
      pp_buf_data_rsci_bcwt_1 <= 1'b0;
    end
    else begin
      pp_buf_data_rsci_bcwt_1 <= ~((~(pp_buf_data_rsci_bcwt_1 | pp_buf_data_rsci_biwt_1))
          | pp_buf_data_rsci_bdwt_2);
    end
  end
  always @(posedge clk) begin
    if ( pp_buf_data_rsci_biwt_1 ) begin
      pp_buf_data_rsci_q_d_bfwt <= pp_buf_data_rsci_q_d;
    end
  end

  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_ctrl
    (
  run_wen, run_wten, pp_buf_data_rsci_oswt_1, pp_buf_data_rsci_biwt_1, pp_buf_data_rsci_bdwt_2,
      pp_buf_data_rsci_we_d_run_sct_pff, pp_buf_data_rsci_iswt0_pff, pp_buf_data_rsci_re_d_run_sct_pff,
      pp_buf_data_rsci_oswt_1_pff
);
  input run_wen;
  input run_wten;
  input pp_buf_data_rsci_oswt_1;
  output pp_buf_data_rsci_biwt_1;
  output pp_buf_data_rsci_bdwt_2;
  output pp_buf_data_rsci_we_d_run_sct_pff;
  input pp_buf_data_rsci_iswt0_pff;
  output pp_buf_data_rsci_re_d_run_sct_pff;
  input pp_buf_data_rsci_oswt_1_pff;



  // Interconnect Declarations for Component Instantiations 
  assign pp_buf_data_rsci_bdwt_2 = pp_buf_data_rsci_oswt_1 & run_wen;
  assign pp_buf_data_rsci_biwt_1 = (~ run_wten) & pp_buf_data_rsci_oswt_1;
  assign pp_buf_data_rsci_we_d_run_sct_pff = pp_buf_data_rsci_iswt0_pff & run_wen;
  assign pp_buf_data_rsci_re_d_run_sct_pff = pp_buf_data_rsci_oswt_1_pff & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_v_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_v_chan1_wait_ctrl (
  v_chan1_rsci_iswt0, v_chan1_rsci_biwt, v_chan1_rsci_irdy
);
  input v_chan1_rsci_iswt0;
  output v_chan1_rsci_biwt;
  input v_chan1_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign v_chan1_rsci_biwt = v_chan1_rsci_iswt0 & v_chan1_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_k_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_k_chan1_wait_ctrl (
  k_chan1_rsci_iswt0, k_chan1_rsci_biwt, k_chan1_rsci_irdy
);
  input k_chan1_rsci_iswt0;
  output k_chan1_rsci_biwt;
  input k_chan1_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign k_chan1_rsci_biwt = k_chan1_rsci_iswt0 & k_chan1_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_q_chan1_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_q_chan1_wait_ctrl (
  q_chan1_rsci_iswt0, q_chan1_rsci_biwt, q_chan1_rsci_irdy
);
  input q_chan1_rsci_iswt0;
  output q_chan1_rsci_biwt;
  input q_chan1_rsci_irdy;



  // Interconnect Declarations for Component Instantiations 
  assign q_chan1_rsci_biwt = q_chan1_rsci_iswt0 & q_chan1_rsci_irdy;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_din_chan_rsci_din_chan_wait_ctrl
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_din_chan_rsci_din_chan_wait_ctrl (
  run_wen, din_chan_rsci_iswt0, din_chan_rsci_irdy_run_sct
);
  input run_wen;
  input din_chan_rsci_iswt0;
  output din_chan_rsci_irdy_run_sct;



  // Interconnect Declarations for Component Instantiations 
  assign din_chan_rsci_irdy_run_sct = din_chan_rsci_iswt0 & run_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1 (
  clk, rst, arst_n, pp_buf_data_rsci_q_d, run_wen, run_wten, pp_buf_data_rsci_oswt_1,
      pp_buf_data_rsci_q_d_mxwt, pp_buf_data_rsci_we_d_pff, pp_buf_data_rsci_iswt0_pff,
      pp_buf_data_rsci_re_d_pff, pp_buf_data_rsci_oswt_1_pff
);
  input clk;
  input rst;
  input arst_n;
  input [15:0] pp_buf_data_rsci_q_d;
  input run_wen;
  input run_wten;
  input pp_buf_data_rsci_oswt_1;
  output [15:0] pp_buf_data_rsci_q_d_mxwt;
  output pp_buf_data_rsci_we_d_pff;
  input pp_buf_data_rsci_iswt0_pff;
  output pp_buf_data_rsci_re_d_pff;
  input pp_buf_data_rsci_oswt_1_pff;


  // Interconnect Declarations
  wire pp_buf_data_rsci_biwt_1;
  wire pp_buf_data_rsci_bdwt_2;
  wire pp_buf_data_rsci_we_d_run_sct_iff;
  wire pp_buf_data_rsci_re_d_run_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_ctrl
      ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .run_wten(run_wten),
      .pp_buf_data_rsci_oswt_1(pp_buf_data_rsci_oswt_1),
      .pp_buf_data_rsci_biwt_1(pp_buf_data_rsci_biwt_1),
      .pp_buf_data_rsci_bdwt_2(pp_buf_data_rsci_bdwt_2),
      .pp_buf_data_rsci_we_d_run_sct_pff(pp_buf_data_rsci_we_d_run_sct_iff),
      .pp_buf_data_rsci_iswt0_pff(pp_buf_data_rsci_iswt0_pff),
      .pp_buf_data_rsci_re_d_run_sct_pff(pp_buf_data_rsci_re_d_run_sct_iff),
      .pp_buf_data_rsci_oswt_1_pff(pp_buf_data_rsci_oswt_1_pff)
    );
  ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_dp ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_pp_buf_data_rsc_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pp_buf_data_rsci_q_d(pp_buf_data_rsci_q_d),
      .pp_buf_data_rsci_q_d_mxwt(pp_buf_data_rsci_q_d_mxwt),
      .pp_buf_data_rsci_biwt_1(pp_buf_data_rsci_biwt_1),
      .pp_buf_data_rsci_bdwt_2(pp_buf_data_rsci_bdwt_2)
    );
  assign pp_buf_data_rsci_we_d_pff = pp_buf_data_rsci_we_d_run_sct_iff;
  assign pp_buf_data_rsci_re_d_pff = pp_buf_data_rsci_re_d_run_sct_iff;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci (
  v_chan1_rsc_dat, v_chan1_rsc_vld, v_chan1_rsc_rdy, v_chan1_rsci_oswt, v_chan1_rsci_wen_comp,
      v_chan1_rsci_idat
);
  output [1023:0] v_chan1_rsc_dat;
  output v_chan1_rsc_vld;
  input v_chan1_rsc_rdy;
  input v_chan1_rsci_oswt;
  output v_chan1_rsci_wen_comp;
  input [1023:0] v_chan1_rsci_idat;


  // Interconnect Declarations
  wire v_chan1_rsci_biwt;
  wire v_chan1_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd7),
  .width(32'sd1024)) v_chan1_rsci (
      .irdy(v_chan1_rsci_irdy),
      .ivld(v_chan1_rsci_oswt),
      .idat(v_chan1_rsci_idat),
      .rdy(v_chan1_rsc_rdy),
      .vld(v_chan1_rsc_vld),
      .dat(v_chan1_rsc_dat)
    );
  ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_v_chan1_wait_ctrl ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_v_chan1_wait_ctrl_inst
      (
      .v_chan1_rsci_iswt0(v_chan1_rsci_oswt),
      .v_chan1_rsci_biwt(v_chan1_rsci_biwt),
      .v_chan1_rsci_irdy(v_chan1_rsci_irdy)
    );
  assign v_chan1_rsci_wen_comp = (~ v_chan1_rsci_oswt) | v_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci (
  k_chan1_rsc_dat, k_chan1_rsc_vld, k_chan1_rsc_rdy, k_chan1_rsci_oswt, k_chan1_rsci_wen_comp,
      k_chan1_rsci_idat
);
  output [1023:0] k_chan1_rsc_dat;
  output k_chan1_rsc_vld;
  input k_chan1_rsc_rdy;
  input k_chan1_rsci_oswt;
  output k_chan1_rsci_wen_comp;
  input [1023:0] k_chan1_rsci_idat;


  // Interconnect Declarations
  wire k_chan1_rsci_biwt;
  wire k_chan1_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd6),
  .width(32'sd1024)) k_chan1_rsci (
      .irdy(k_chan1_rsci_irdy),
      .ivld(k_chan1_rsci_oswt),
      .idat(k_chan1_rsci_idat),
      .rdy(k_chan1_rsc_rdy),
      .vld(k_chan1_rsc_vld),
      .dat(k_chan1_rsc_dat)
    );
  ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_k_chan1_wait_ctrl ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_k_chan1_wait_ctrl_inst
      (
      .k_chan1_rsci_iswt0(k_chan1_rsci_oswt),
      .k_chan1_rsci_biwt(k_chan1_rsci_biwt),
      .k_chan1_rsci_irdy(k_chan1_rsci_irdy)
    );
  assign k_chan1_rsci_wen_comp = (~ k_chan1_rsci_oswt) | k_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci (
  q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy, q_chan1_rsci_oswt, q_chan1_rsci_wen_comp,
      q_chan1_rsci_idat
);
  output [1023:0] q_chan1_rsc_dat;
  output q_chan1_rsc_vld;
  input q_chan1_rsc_rdy;
  input q_chan1_rsci_oswt;
  output q_chan1_rsci_wen_comp;
  input [1023:0] q_chan1_rsci_idat;


  // Interconnect Declarations
  wire q_chan1_rsci_biwt;
  wire q_chan1_rsci_irdy;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd5),
  .width(32'sd1024)) q_chan1_rsci (
      .irdy(q_chan1_rsci_irdy),
      .ivld(q_chan1_rsci_oswt),
      .idat(q_chan1_rsci_idat),
      .rdy(q_chan1_rsc_rdy),
      .vld(q_chan1_rsc_vld),
      .dat(q_chan1_rsc_dat)
    );
  ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_q_chan1_wait_ctrl ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_q_chan1_wait_ctrl_inst
      (
      .q_chan1_rsci_iswt0(q_chan1_rsci_oswt),
      .q_chan1_rsci_biwt(q_chan1_rsci_biwt),
      .q_chan1_rsci_irdy(q_chan1_rsci_irdy)
    );
  assign q_chan1_rsci_wen_comp = (~ q_chan1_rsci_oswt) | q_chan1_rsci_biwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run_din_chan_rsci
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run_din_chan_rsci (
  din_chan_rsc_dat, din_chan_rsc_vld, din_chan_rsc_rdy, run_wen, din_chan_rsci_oswt,
      din_chan_rsci_wen_comp, din_chan_rsci_idat_mxwt
);
  input [15:0] din_chan_rsc_dat;
  input din_chan_rsc_vld;
  output din_chan_rsc_rdy;
  input run_wen;
  input din_chan_rsci_oswt;
  output din_chan_rsci_wen_comp;
  output [15:0] din_chan_rsci_idat_mxwt;


  // Interconnect Declarations
  wire din_chan_rsci_irdy_run_sct;
  wire din_chan_rsci_ivld;
  wire [15:0] din_chan_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_coupled_v1 #(.rscid(32'sd4),
  .width(32'sd16)) din_chan_rsci (
      .rdy(din_chan_rsc_rdy),
      .vld(din_chan_rsc_vld),
      .dat(din_chan_rsc_dat),
      .irdy(din_chan_rsci_irdy_run_sct),
      .ivld(din_chan_rsci_ivld),
      .idat(din_chan_rsci_idat)
    );
  ATTENTION_IP_Attention_Buffer_run_din_chan_rsci_din_chan_wait_ctrl ATTENTION_IP_Attention_Buffer_run_din_chan_rsci_din_chan_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .din_chan_rsci_iswt0(din_chan_rsci_oswt),
      .din_chan_rsci_irdy_run_sct(din_chan_rsci_irdy_run_sct)
    );
  assign din_chan_rsci_idat_mxwt = din_chan_rsci_idat;
  assign din_chan_rsci_wen_comp = (~ din_chan_rsci_oswt) | din_chan_rsci_ivld;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer_run
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer_run (
  clk, rst, arst_n, head, length, dim, din_chan_rsc_dat, din_chan_rsc_vld, din_chan_rsc_rdy,
      q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy, k_chan1_rsc_dat, k_chan1_rsc_vld,
      k_chan1_rsc_rdy, v_chan1_rsc_dat, v_chan1_rsc_vld, v_chan1_rsc_rdy, pp_buf_data_rsci_radr_d,
      pp_buf_data_rsci_wadr_d, pp_buf_data_rsci_d_d, pp_buf_data_rsci_q_d, pp_buf_data_rsci_we_d_pff,
      pp_buf_data_rsci_re_d_pff
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [15:0] din_chan_rsc_dat;
  input din_chan_rsc_vld;
  output din_chan_rsc_rdy;
  output [1023:0] q_chan1_rsc_dat;
  output q_chan1_rsc_vld;
  input q_chan1_rsc_rdy;
  output [1023:0] k_chan1_rsc_dat;
  output k_chan1_rsc_vld;
  input k_chan1_rsc_rdy;
  output [1023:0] v_chan1_rsc_dat;
  output v_chan1_rsc_vld;
  input v_chan1_rsc_rdy;
  output [13:0] pp_buf_data_rsci_radr_d;
  output [13:0] pp_buf_data_rsci_wadr_d;
  output [15:0] pp_buf_data_rsci_d_d;
  input [15:0] pp_buf_data_rsci_q_d;
  output pp_buf_data_rsci_we_d_pff;
  output pp_buf_data_rsci_re_d_pff;


  // Interconnect Declarations
  wire run_wen;
  wire run_wten;
  wire din_chan_rsci_wen_comp;
  wire [15:0] din_chan_rsci_idat_mxwt;
  wire q_chan1_rsci_wen_comp;
  wire k_chan1_rsci_wen_comp;
  wire v_chan1_rsci_wen_comp;
  wire [15:0] pp_buf_data_rsci_q_d_mxwt;
  reg [15:0] q_chan1_rsci_idat_1023_1008;
  reg [15:0] q_chan1_rsci_idat_1007_992;
  reg [15:0] q_chan1_rsci_idat_991_976;
  reg [15:0] q_chan1_rsci_idat_975_960;
  reg [15:0] q_chan1_rsci_idat_959_944;
  reg [15:0] q_chan1_rsci_idat_943_928;
  reg [15:0] q_chan1_rsci_idat_927_912;
  reg [15:0] q_chan1_rsci_idat_911_896;
  reg [15:0] q_chan1_rsci_idat_895_880;
  reg [15:0] q_chan1_rsci_idat_879_864;
  reg [15:0] q_chan1_rsci_idat_863_848;
  reg [15:0] q_chan1_rsci_idat_847_832;
  reg [15:0] q_chan1_rsci_idat_831_816;
  reg [15:0] q_chan1_rsci_idat_815_800;
  reg [15:0] q_chan1_rsci_idat_799_784;
  reg [15:0] q_chan1_rsci_idat_783_768;
  reg [15:0] q_chan1_rsci_idat_767_752;
  reg [15:0] q_chan1_rsci_idat_751_736;
  reg [15:0] q_chan1_rsci_idat_735_720;
  reg [15:0] q_chan1_rsci_idat_719_704;
  reg [15:0] q_chan1_rsci_idat_703_688;
  reg [15:0] q_chan1_rsci_idat_687_672;
  reg [15:0] q_chan1_rsci_idat_671_656;
  reg [15:0] q_chan1_rsci_idat_655_640;
  reg [15:0] q_chan1_rsci_idat_639_624;
  reg [15:0] q_chan1_rsci_idat_623_608;
  reg [15:0] q_chan1_rsci_idat_607_592;
  reg [15:0] q_chan1_rsci_idat_591_576;
  reg [15:0] q_chan1_rsci_idat_575_560;
  reg [15:0] q_chan1_rsci_idat_559_544;
  reg [15:0] q_chan1_rsci_idat_543_528;
  reg [15:0] q_chan1_rsci_idat_527_512;
  reg [15:0] q_chan1_rsci_idat_511_496;
  reg [15:0] q_chan1_rsci_idat_495_480;
  reg [15:0] q_chan1_rsci_idat_479_464;
  reg [15:0] q_chan1_rsci_idat_463_448;
  reg [15:0] q_chan1_rsci_idat_447_432;
  reg [15:0] q_chan1_rsci_idat_431_416;
  reg [15:0] q_chan1_rsci_idat_415_400;
  reg [15:0] q_chan1_rsci_idat_399_384;
  reg [15:0] q_chan1_rsci_idat_383_368;
  reg [15:0] q_chan1_rsci_idat_367_352;
  reg [15:0] q_chan1_rsci_idat_351_336;
  reg [15:0] q_chan1_rsci_idat_335_320;
  reg [15:0] q_chan1_rsci_idat_319_304;
  reg [15:0] q_chan1_rsci_idat_303_288;
  reg [15:0] q_chan1_rsci_idat_287_272;
  reg [15:0] q_chan1_rsci_idat_271_256;
  reg [15:0] q_chan1_rsci_idat_255_240;
  reg [15:0] q_chan1_rsci_idat_239_224;
  reg [15:0] q_chan1_rsci_idat_223_208;
  reg [15:0] q_chan1_rsci_idat_207_192;
  reg [15:0] q_chan1_rsci_idat_191_176;
  reg [15:0] q_chan1_rsci_idat_175_160;
  reg [15:0] q_chan1_rsci_idat_159_144;
  reg [15:0] q_chan1_rsci_idat_143_128;
  reg [15:0] q_chan1_rsci_idat_127_112;
  reg [15:0] q_chan1_rsci_idat_111_96;
  reg [15:0] q_chan1_rsci_idat_95_80;
  reg [15:0] q_chan1_rsci_idat_79_64;
  reg [15:0] q_chan1_rsci_idat_63_48;
  reg [15:0] q_chan1_rsci_idat_47_32;
  reg [15:0] q_chan1_rsci_idat_31_16;
  reg [15:0] q_chan1_rsci_idat_15_0;
  reg [15:0] k_chan1_rsci_idat_1023_1008;
  reg [15:0] k_chan1_rsci_idat_1007_992;
  reg [15:0] k_chan1_rsci_idat_991_976;
  reg [15:0] k_chan1_rsci_idat_975_960;
  reg [15:0] k_chan1_rsci_idat_959_944;
  reg [15:0] k_chan1_rsci_idat_943_928;
  reg [15:0] k_chan1_rsci_idat_927_912;
  reg [15:0] k_chan1_rsci_idat_911_896;
  reg [15:0] k_chan1_rsci_idat_895_880;
  reg [15:0] k_chan1_rsci_idat_879_864;
  reg [15:0] k_chan1_rsci_idat_863_848;
  reg [15:0] k_chan1_rsci_idat_847_832;
  reg [15:0] k_chan1_rsci_idat_831_816;
  reg [15:0] k_chan1_rsci_idat_815_800;
  reg [15:0] k_chan1_rsci_idat_799_784;
  reg [15:0] k_chan1_rsci_idat_783_768;
  reg [15:0] k_chan1_rsci_idat_767_752;
  reg [15:0] k_chan1_rsci_idat_751_736;
  reg [15:0] k_chan1_rsci_idat_735_720;
  reg [15:0] k_chan1_rsci_idat_719_704;
  reg [15:0] k_chan1_rsci_idat_703_688;
  reg [15:0] k_chan1_rsci_idat_687_672;
  reg [15:0] k_chan1_rsci_idat_671_656;
  reg [15:0] k_chan1_rsci_idat_655_640;
  reg [15:0] k_chan1_rsci_idat_639_624;
  reg [15:0] k_chan1_rsci_idat_623_608;
  reg [15:0] k_chan1_rsci_idat_607_592;
  reg [15:0] k_chan1_rsci_idat_591_576;
  reg [15:0] k_chan1_rsci_idat_575_560;
  reg [15:0] k_chan1_rsci_idat_559_544;
  reg [15:0] k_chan1_rsci_idat_543_528;
  reg [15:0] k_chan1_rsci_idat_527_512;
  reg [15:0] k_chan1_rsci_idat_511_496;
  reg [15:0] k_chan1_rsci_idat_495_480;
  reg [15:0] k_chan1_rsci_idat_479_464;
  reg [15:0] k_chan1_rsci_idat_463_448;
  reg [15:0] k_chan1_rsci_idat_447_432;
  reg [15:0] k_chan1_rsci_idat_431_416;
  reg [15:0] k_chan1_rsci_idat_415_400;
  reg [15:0] k_chan1_rsci_idat_399_384;
  reg [15:0] k_chan1_rsci_idat_383_368;
  reg [15:0] k_chan1_rsci_idat_367_352;
  reg [15:0] k_chan1_rsci_idat_351_336;
  reg [15:0] k_chan1_rsci_idat_335_320;
  reg [15:0] k_chan1_rsci_idat_319_304;
  reg [15:0] k_chan1_rsci_idat_303_288;
  reg [15:0] k_chan1_rsci_idat_287_272;
  reg [15:0] k_chan1_rsci_idat_271_256;
  reg [15:0] k_chan1_rsci_idat_255_240;
  reg [15:0] k_chan1_rsci_idat_239_224;
  reg [15:0] k_chan1_rsci_idat_223_208;
  reg [15:0] k_chan1_rsci_idat_207_192;
  reg [15:0] k_chan1_rsci_idat_191_176;
  reg [15:0] k_chan1_rsci_idat_175_160;
  reg [15:0] k_chan1_rsci_idat_159_144;
  reg [15:0] k_chan1_rsci_idat_143_128;
  reg [15:0] k_chan1_rsci_idat_127_112;
  reg [15:0] k_chan1_rsci_idat_111_96;
  reg [15:0] k_chan1_rsci_idat_95_80;
  reg [15:0] k_chan1_rsci_idat_79_64;
  reg [15:0] k_chan1_rsci_idat_63_48;
  reg [15:0] k_chan1_rsci_idat_47_32;
  reg [15:0] k_chan1_rsci_idat_31_16;
  reg [15:0] k_chan1_rsci_idat_15_0;
  reg [15:0] v_chan1_rsci_idat_1023_1008;
  reg [15:0] v_chan1_rsci_idat_1007_992;
  reg [15:0] v_chan1_rsci_idat_991_976;
  reg [15:0] v_chan1_rsci_idat_975_960;
  reg [15:0] v_chan1_rsci_idat_959_944;
  reg [15:0] v_chan1_rsci_idat_943_928;
  reg [15:0] v_chan1_rsci_idat_927_912;
  reg [15:0] v_chan1_rsci_idat_911_896;
  reg [15:0] v_chan1_rsci_idat_895_880;
  reg [15:0] v_chan1_rsci_idat_879_864;
  reg [15:0] v_chan1_rsci_idat_863_848;
  reg [15:0] v_chan1_rsci_idat_847_832;
  reg [15:0] v_chan1_rsci_idat_831_816;
  reg [15:0] v_chan1_rsci_idat_815_800;
  reg [15:0] v_chan1_rsci_idat_799_784;
  reg [15:0] v_chan1_rsci_idat_783_768;
  reg [15:0] v_chan1_rsci_idat_767_752;
  reg [15:0] v_chan1_rsci_idat_751_736;
  reg [15:0] v_chan1_rsci_idat_735_720;
  reg [15:0] v_chan1_rsci_idat_719_704;
  reg [15:0] v_chan1_rsci_idat_703_688;
  reg [15:0] v_chan1_rsci_idat_687_672;
  reg [15:0] v_chan1_rsci_idat_671_656;
  reg [15:0] v_chan1_rsci_idat_655_640;
  reg [15:0] v_chan1_rsci_idat_639_624;
  reg [15:0] v_chan1_rsci_idat_623_608;
  reg [15:0] v_chan1_rsci_idat_607_592;
  reg [15:0] v_chan1_rsci_idat_591_576;
  reg [15:0] v_chan1_rsci_idat_575_560;
  reg [15:0] v_chan1_rsci_idat_559_544;
  reg [15:0] v_chan1_rsci_idat_543_528;
  reg [15:0] v_chan1_rsci_idat_527_512;
  reg [15:0] v_chan1_rsci_idat_511_496;
  reg [15:0] v_chan1_rsci_idat_495_480;
  reg [15:0] v_chan1_rsci_idat_479_464;
  reg [15:0] v_chan1_rsci_idat_463_448;
  reg [15:0] v_chan1_rsci_idat_447_432;
  reg [15:0] v_chan1_rsci_idat_431_416;
  reg [15:0] v_chan1_rsci_idat_415_400;
  reg [15:0] v_chan1_rsci_idat_399_384;
  reg [15:0] v_chan1_rsci_idat_383_368;
  reg [15:0] v_chan1_rsci_idat_367_352;
  reg [15:0] v_chan1_rsci_idat_351_336;
  reg [15:0] v_chan1_rsci_idat_335_320;
  reg [15:0] v_chan1_rsci_idat_319_304;
  reg [15:0] v_chan1_rsci_idat_303_288;
  reg [15:0] v_chan1_rsci_idat_287_272;
  reg [15:0] v_chan1_rsci_idat_271_256;
  reg [15:0] v_chan1_rsci_idat_255_240;
  reg [15:0] v_chan1_rsci_idat_239_224;
  reg [15:0] v_chan1_rsci_idat_223_208;
  reg [15:0] v_chan1_rsci_idat_207_192;
  reg [15:0] v_chan1_rsci_idat_191_176;
  reg [15:0] v_chan1_rsci_idat_175_160;
  reg [15:0] v_chan1_rsci_idat_159_144;
  reg [15:0] v_chan1_rsci_idat_143_128;
  reg [15:0] v_chan1_rsci_idat_127_112;
  reg [15:0] v_chan1_rsci_idat_111_96;
  reg [15:0] v_chan1_rsci_idat_95_80;
  reg [15:0] v_chan1_rsci_idat_79_64;
  reg [15:0] v_chan1_rsci_idat_63_48;
  reg [15:0] v_chan1_rsci_idat_47_32;
  reg [15:0] v_chan1_rsci_idat_31_16;
  reg [15:0] v_chan1_rsci_idat_15_0;
  wire [8:0] fsm_output;
  wire LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp;
  wire LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp;
  wire LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp;
  wire [6:0] LOOPK1_acc_1_tmp;
  wire [7:0] nl_LOOPK1_acc_1_tmp;
  wire or_dcpl;
  wire or_dcpl_1;
  wire or_dcpl_2;
  wire or_dcpl_3;
  wire or_dcpl_4;
  wire or_dcpl_6;
  wire or_dcpl_8;
  wire or_dcpl_9;
  wire or_dcpl_10;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire or_dcpl_14;
  wire or_dcpl_15;
  wire or_dcpl_17;
  wire or_dcpl_18;
  wire or_dcpl_20;
  wire or_dcpl_22;
  wire or_dcpl_30;
  wire or_dcpl_33;
  wire or_dcpl_34;
  wire or_dcpl_36;
  wire or_dcpl_37;
  wire or_dcpl_53;
  wire or_dcpl_55;
  wire or_dcpl_71;
  wire or_dcpl_73;
  wire and_dcpl_7;
  wire and_dcpl_8;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_12;
  wire and_dcpl_14;
  wire and_dcpl_15;
  wire and_dcpl_16;
  wire and_dcpl_18;
  wire or_dcpl_93;
  wire or_dcpl_99;
  wire or_dcpl_101;
  wire or_dcpl_104;
  wire or_dcpl_109;
  wire or_dcpl_113;
  wire or_dcpl_114;
  wire and_dcpl_23;
  wire and_dcpl_24;
  wire or_tmp_23;
  wire mux_tmp_26;
  wire mux_tmp_27;
  wire mux_tmp_31;
  wire mux_tmp_34;
  wire and_dcpl_32;
  wire and_dcpl_33;
  wire and_dcpl_34;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire and_dcpl_38;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire or_dcpl_121;
  wire or_dcpl_122;
  wire or_dcpl_123;
  wire or_dcpl_124;
  wire or_dcpl_126;
  wire or_dcpl_127;
  wire or_dcpl_129;
  wire or_dcpl_130;
  wire or_dcpl_131;
  wire or_dcpl_132;
  wire or_dcpl_134;
  wire or_dcpl_136;
  wire or_dcpl_138;
  wire or_dcpl_139;
  wire or_dcpl_141;
  wire or_dcpl_149;
  wire or_dcpl_152;
  wire or_dcpl_153;
  wire or_dcpl_155;
  wire or_dcpl_156;
  wire or_dcpl_172;
  wire or_dcpl_174;
  wire or_dcpl_190;
  wire or_dcpl_192;
  wire or_tmp_46;
  wire mux_tmp_53;
  wire mux_tmp_58;
  wire mux_tmp_59;
  wire mux_tmp_62;
  wire or_tmp_51;
  wire or_tmp_53;
  wire and_dcpl_51;
  wire mux_tmp_74;
  wire and_dcpl_53;
  wire mux_tmp_83;
  wire and_dcpl_54;
  wire and_dcpl_55;
  wire nor_tmp_13;
  wire or_tmp_70;
  wire mux_tmp_90;
  wire mux_tmp_91;
  wire and_dcpl_57;
  wire or_tmp_74;
  wire mux_tmp_92;
  wire mux_tmp_93;
  wire mux_tmp_94;
  wire mux_tmp_95;
  wire and_dcpl_61;
  wire and_dcpl_63;
  wire mux_tmp_96;
  wire and_dcpl_65;
  wire and_dcpl_68;
  wire and_dcpl_69;
  wire mux_tmp_97;
  wire and_dcpl_71;
  wire and_dcpl_72;
  wire mux_tmp_98;
  wire and_dcpl_76;
  wire and_dcpl_77;
  wire and_dcpl_79;
  wire and_dcpl_83;
  wire and_dcpl_84;
  wire and_dcpl_86;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_93;
  wire mux_tmp_99;
  wire mux_tmp_100;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_104;
  wire and_dcpl_105;
  wire and_dcpl_109;
  wire and_dcpl_111;
  wire and_dcpl_115;
  wire and_dcpl_117;
  wire and_dcpl_121;
  wire and_dcpl_123;
  wire and_dcpl_127;
  wire and_dcpl_129;
  wire and_dcpl_133;
  wire and_dcpl_135;
  wire and_dcpl_139;
  wire and_dcpl_141;
  wire mux_tmp_102;
  wire or_tmp_96;
  wire mux_tmp_104;
  wire mux_tmp_105;
  wire mux_tmp_106;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire and_dcpl_155;
  wire and_dcpl_156;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire and_dcpl_163;
  wire and_dcpl_164;
  wire and_dcpl_165;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_168;
  wire and_dcpl_169;
  wire and_dcpl_170;
  wire and_dcpl_171;
  wire and_dcpl_172;
  wire and_dcpl_173;
  wire and_dcpl_174;
  wire and_dcpl_175;
  wire and_dcpl_176;
  wire and_dcpl_177;
  wire and_dcpl_178;
  wire and_dcpl_179;
  wire and_dcpl_180;
  wire and_dcpl_181;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_195;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire and_dcpl_201;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_204;
  wire and_dcpl_205;
  wire and_dcpl_206;
  wire and_dcpl_207;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire and_dcpl_213;
  wire and_dcpl_214;
  wire and_dcpl_215;
  wire and_dcpl_216;
  wire and_dcpl_217;
  wire and_dcpl_218;
  wire or_dcpl_219;
  wire or_dcpl_220;
  wire or_dcpl_222;
  wire or_dcpl_226;
  wire or_dcpl_227;
  wire or_dcpl_228;
  wire or_dcpl_230;
  wire or_dcpl_232;
  wire or_dcpl_235;
  wire or_dcpl_236;
  wire or_dcpl_238;
  wire or_dcpl_239;
  wire or_dcpl_243;
  wire or_dcpl_244;
  wire or_dcpl_246;
  wire or_dcpl_250;
  wire or_dcpl_251;
  wire or_dcpl_253;
  wire or_dcpl_257;
  wire or_dcpl_258;
  wire or_dcpl_260;
  wire or_dcpl_268;
  wire or_dcpl_269;
  wire or_dcpl_271;
  wire or_dcpl_272;
  wire or_dcpl_276;
  wire or_dcpl_278;
  wire or_dcpl_282;
  wire or_dcpl_284;
  wire or_dcpl_288;
  wire or_dcpl_290;
  wire or_dcpl_294;
  wire or_dcpl_296;
  wire or_dcpl_300;
  wire or_dcpl_302;
  wire or_dcpl_306;
  wire or_dcpl_308;
  wire mux_tmp_140;
  wire mux_tmp_143;
  reg LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm;
  wire LOOPK3_and_cse;
  wire LOOPK2_and_cse;
  wire LOOPJ2_and_cse;
  wire channel_in_data_and_cse;
  reg reg_din_chan_rsci_oswt_cse;
  reg reg_q_chan1_rsci_oswt_cse;
  reg reg_k_chan1_rsci_oswt_cse;
  reg reg_v_chan1_rsci_oswt_cse;
  reg reg_pp_buf_data_rsci_oswt_1_cse;
  wire or_108_cse;
  wire and_237_cse;
  wire nor_49_cse;
  wire or_145_cse;
  wire or_111_cse;
  wire nor_28_cse;
  wire or_319_cse;
  wire nor_34_cse;
  wire [7:0] LOOPJ1_acc_sdt;
  wire [8:0] nl_LOOPJ1_acc_sdt;
  reg LOOPJ1_acc_itm_7;
  reg [6:0] LOOPJ1_acc_itm_6_0;
  wire LOOPJ1_j_and_ssc;
  wire nor_53_cse;
  wire nor_54_cse;
  wire mux_16_cse;
  wire pp_buf_data_rsci_we_d_iff;
  wire pp_buf_data_rsci_re_d_iff;
  reg [15:0] channel_in_data_63_lpi_4;
  reg [15:0] LOOPJ2_asn_itm;
  reg [15:0] channel_in_data_62_lpi_4;
  reg [15:0] channel_in_data_1_lpi_4;
  reg [15:0] channel_in_data_61_lpi_4;
  reg [15:0] channel_in_data_2_lpi_4;
  reg [15:0] channel_in_data_60_lpi_4;
  reg [15:0] channel_in_data_3_lpi_4;
  reg [15:0] channel_in_data_59_lpi_4;
  reg [15:0] channel_in_data_4_lpi_4;
  reg [15:0] channel_in_data_58_lpi_4;
  reg [15:0] channel_in_data_5_lpi_4;
  reg [15:0] channel_in_data_57_lpi_4;
  reg [15:0] channel_in_data_6_lpi_4;
  reg [15:0] channel_in_data_56_lpi_4;
  reg [15:0] channel_in_data_7_lpi_4;
  reg [15:0] channel_in_data_55_lpi_4;
  reg [15:0] channel_in_data_8_lpi_4;
  reg [15:0] channel_in_data_54_lpi_4;
  reg [15:0] channel_in_data_9_lpi_4;
  reg [15:0] channel_in_data_53_lpi_4;
  reg [15:0] channel_in_data_10_lpi_4;
  reg [15:0] channel_in_data_52_lpi_4;
  reg [15:0] channel_in_data_11_lpi_4;
  reg [15:0] channel_in_data_51_lpi_4;
  reg [15:0] channel_in_data_12_lpi_4;
  reg [15:0] channel_in_data_50_lpi_4;
  reg [15:0] channel_in_data_13_lpi_4;
  reg [15:0] channel_in_data_49_lpi_4;
  reg [15:0] channel_in_data_14_lpi_4;
  reg [15:0] channel_in_data_48_lpi_4;
  reg [15:0] channel_in_data_15_lpi_4;
  reg [15:0] channel_in_data_47_lpi_4;
  reg [15:0] channel_in_data_16_lpi_4;
  reg [15:0] channel_in_data_46_lpi_4;
  reg [15:0] channel_in_data_17_lpi_4;
  reg [15:0] channel_in_data_45_lpi_4;
  reg [15:0] channel_in_data_18_lpi_4;
  reg [15:0] channel_in_data_44_lpi_4;
  reg [15:0] channel_in_data_19_lpi_4;
  reg [15:0] channel_in_data_43_lpi_4;
  reg [15:0] channel_in_data_20_lpi_4;
  reg [15:0] channel_in_data_42_lpi_4;
  reg [15:0] channel_in_data_21_lpi_4;
  reg [15:0] channel_in_data_41_lpi_4;
  reg [15:0] channel_in_data_22_lpi_4;
  reg [15:0] channel_in_data_40_lpi_4;
  reg [15:0] channel_in_data_23_lpi_4;
  reg [15:0] channel_in_data_39_lpi_4;
  reg [15:0] channel_in_data_24_lpi_4;
  reg [15:0] channel_in_data_38_lpi_4;
  reg [15:0] channel_in_data_25_lpi_4;
  reg [15:0] channel_in_data_37_lpi_4;
  reg [15:0] channel_in_data_26_lpi_4;
  reg [15:0] channel_in_data_36_lpi_4;
  reg [15:0] channel_in_data_27_lpi_4;
  reg [15:0] channel_in_data_35_lpi_4;
  reg [15:0] channel_in_data_28_lpi_4;
  reg [15:0] channel_in_data_34_lpi_4;
  reg [15:0] channel_in_data_29_lpi_4;
  reg [15:0] channel_in_data_33_lpi_4;
  reg [15:0] channel_in_data_30_lpi_4;
  reg [15:0] channel_in_data_32_lpi_4;
  reg [15:0] channel_in_data_31_lpi_4;
  reg [5:0] LOOPJ1_j_sva_5_0;
  wire [6:0] LOOPK2_acc_tmp_sva_mx0w2;
  wire [7:0] nl_LOOPK2_acc_tmp_sva_mx0w2;
  reg [5:0] LOOPK2_acc_1_itm;
  wire [6:0] LOOPK3_acc_psp_sva_mx0w4;
  wire [7:0] nl_LOOPK3_acc_psp_sva_mx0w4;
  reg LOOPJ1_j_sva_7;
  reg LOOPJ1_j_sva_6;
  wire mux_69_itm;
  wire mux_110_itm;
  wire and_dcpl;
  wire and_dcpl_227;
  wire [5:0] z_out;
  wire [6:0] nl_z_out;
  wire and_dcpl_246;
  wire [7:0] z_out_1;
  wire [8:0] nl_z_out_1;
  reg [3:0] LOOPI1_i_sva;
  reg [5:0] LOOPK3_acc_1_itm;
  reg [15:0] LOOPJ2_asn_itm_1;
  reg [15:0] LOOPJ2_asn_itm_2;
  reg [15:0] LOOPJ2_asn_itm_3;
  reg [15:0] LOOPJ2_asn_itm_4;
  reg [15:0] LOOPJ2_asn_itm_5;
  reg [15:0] LOOPJ2_asn_itm_6;
  reg [15:0] LOOPJ2_asn_itm_7;
  reg [15:0] LOOPJ2_asn_itm_8;
  reg [15:0] LOOPJ2_asn_itm_9;
  reg [15:0] LOOPJ2_asn_itm_10;
  reg [15:0] LOOPJ2_asn_itm_11;
  reg [15:0] LOOPJ2_asn_itm_12;
  reg [15:0] LOOPJ2_asn_itm_13;
  reg [15:0] LOOPJ2_asn_itm_14;
  reg [15:0] LOOPJ2_asn_itm_15;
  reg [15:0] LOOPJ2_asn_itm_16;
  reg [15:0] LOOPJ2_asn_itm_17;
  reg [15:0] LOOPJ2_asn_itm_18;
  reg [15:0] LOOPJ2_asn_itm_19;
  reg [15:0] LOOPJ2_asn_itm_20;
  reg [15:0] LOOPJ2_asn_itm_21;
  reg [15:0] LOOPJ2_asn_itm_22;
  reg [15:0] LOOPJ2_asn_itm_23;
  reg [15:0] LOOPJ2_asn_itm_24;
  reg [15:0] LOOPJ2_asn_itm_25;
  reg [15:0] LOOPJ2_asn_itm_26;
  reg [15:0] LOOPJ2_asn_itm_27;
  reg [15:0] LOOPJ2_asn_itm_28;
  reg [15:0] LOOPJ2_asn_itm_29;
  reg [15:0] LOOPJ2_asn_itm_30;
  reg [15:0] LOOPJ2_asn_itm_31;
  reg [15:0] LOOPJ2_asn_itm_32;
  reg [15:0] LOOPJ2_asn_itm_33;
  reg [15:0] LOOPJ2_asn_itm_34;
  reg [15:0] LOOPJ2_asn_itm_35;
  reg [15:0] LOOPJ2_asn_itm_36;
  reg [15:0] LOOPJ2_asn_itm_37;
  reg [15:0] LOOPJ2_asn_itm_38;
  reg [15:0] LOOPJ2_asn_itm_39;
  reg [15:0] LOOPJ2_asn_itm_40;
  reg [15:0] LOOPJ2_asn_itm_41;
  reg [15:0] LOOPJ2_asn_itm_42;
  reg [15:0] LOOPJ2_asn_itm_43;
  reg [15:0] LOOPJ2_asn_itm_44;
  reg [15:0] LOOPJ2_asn_itm_45;
  reg [15:0] LOOPJ2_asn_itm_46;
  reg [15:0] LOOPJ2_asn_itm_47;
  reg [15:0] LOOPJ2_asn_itm_48;
  reg [15:0] LOOPJ2_asn_itm_49;
  reg [15:0] LOOPJ2_asn_itm_50;
  reg [15:0] LOOPJ2_asn_itm_51;
  reg [15:0] LOOPJ2_asn_itm_52;
  reg [15:0] LOOPJ2_asn_itm_53;
  reg [15:0] LOOPJ2_asn_itm_54;
  reg [15:0] LOOPJ2_asn_itm_55;
  reg [15:0] LOOPJ2_asn_itm_56;
  reg [15:0] LOOPJ2_asn_itm_57;
  reg [15:0] LOOPJ2_asn_itm_58;
  reg [15:0] LOOPJ2_asn_itm_59;
  reg [15:0] LOOPJ2_asn_itm_60;
  reg [15:0] LOOPJ2_asn_itm_61;
  reg [15:0] LOOPJ2_asn_itm_62;
  wire LOOPI1_i_sva_mx0c0;
  wire LOOPJ1_j_sva_mx0c2;
  wire [8:0] operator_6_false_acc_psp_sva_1;
  wire [9:0] nl_operator_6_false_acc_psp_sva_1;
  wire or_146_cse_1;
  wire or_158_cse_1;
  wire or_478_cse;
  wire or_472_cse;
  wire or_476_cse;
  wire nor_145_cse;
  wire mux_36_itm;
  wire and_252_itm;
  wire and_263_itm;
  wire and_271_itm;
  wire and_277_itm;
  wire and_280_itm;
  wire and_286_itm;
  wire nor_63_cse;

  wire LOOPI1_i_not_1_nl;
  wire mux_57_nl;
  wire mux_56_nl;
  wire mux_55_nl;
  wire mux_54_nl;
  wire or_259_nl;
  wire mux_52_nl;
  wire mux_51_nl;
  wire or_258_nl;
  wire or_255_nl;
  wire or_254_nl;
  wire mux_68_nl;
  wire mux_67_nl;
  wire mux_66_nl;
  wire mux_65_nl;
  wire mux_64_nl;
  wire mux_63_nl;
  wire mux_60_nl;
  wire[5:0] LOOPJ2_j_LOOPJ2_j_mux_nl;
  wire and_223_nl;
  wire LOOPK2_not_nl;
  wire mux_148_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire mux_145_nl;
  wire mux_144_nl;
  wire or_452_nl;
  wire mux_142_nl;
  wire or_451_nl;
  wire mux_141_nl;
  wire or_450_nl;
  wire mux_162_nl;
  wire mux_161_nl;
  wire mux_160_nl;
  wire mux_159_nl;
  wire or_475_nl;
  wire mux_158_nl;
  wire mux_nl;
  wire nor_135_nl;
  wire or_473_nl;
  wire mux_155_nl;
  wire or_143_nl;
  wire mux_30_nl;
  wire mux_29_nl;
  wire mux_33_nl;
  wire mux_32_nl;
  wire mux_61_nl;
  wire mux_73_nl;
  wire mux_72_nl;
  wire mux_71_nl;
  wire or_268_nl;
  wire mux_70_nl;
  wire mux_80_nl;
  wire mux_79_nl;
  wire mux_78_nl;
  wire mux_77_nl;
  wire mux_76_nl;
  wire mux_75_nl;
  wire or_270_nl;
  wire or_286_nl;
  wire or_283_nl;
  wire or_287_nl;
  wire nand_12_nl;
  wire nand_nl;
  wire or_292_nl;
  wire nand_14_nl;
  wire or_293_nl;
  wire nand_1_nl;
  wire or_297_nl;
  wire nand_16_nl;
  wire or_299_nl;
  wire or_305_nl;
  wire nand_2_nl;
  wire mux_101_nl;
  wire nor_40_nl;
  wire nor_41_nl;
  wire or_311_nl;
  wire mux_103_nl;
  wire or_309_nl;
  wire nand_17_nl;
  wire mux_107_nl;
  wire nand_18_nl;
  wire or_453_nl;
  wire mux_35_nl;
  wire or_141_nl;
  wire mux_25_nl;
  wire nor_33_nl;
  wire and_nl;
  wire mux_109_nl;
  wire mux_108_nl;
  wire or_105_nl;
  wire[5:0] LOOPJ1_mux_65_nl;
  wire nor_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_165_nl;
  wire mux_164_nl;
  wire nor_136_nl;
  wire nor_137_nl;
  wire nor_138_nl;
  wire mux_163_nl;
  wire nand_27_nl;
  wire or_479_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire mux_123_nl;
  wire mux_122_nl;
  wire mux_121_nl;
  wire nor_55_nl;
  wire or_346_nl;
  wire mux_129_nl;
  wire or_344_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire mux_126_nl;
  wire or_340_nl;
  wire or_326_nl;
  wire[6:0] LOOPK1_k_and_nl;
  wire[6:0] LOOPK1_k_mux1h_nl;
  wire mux_45_nl;
  wire mux_44_nl;
  wire nor_59_nl;
  wire mux_43_nl;
  wire or_466_nl;
  wire or_467_nl;
  wire nor_60_nl;
  wire mux_169_nl;
  wire mux_168_nl;
  wire nor_141_nl;
  wire nor_142_nl;
  wire mux_167_nl;
  wire nor_143_nl;
  wire mux_166_nl;
  wire or_487_nl;
  wire or_486_nl;
  wire nor_144_nl;
  wire LOOPJ1_LOOPJ1_and_nl;
  wire LOOPJ1_mux_nl;
  wire LOOPJ1_and_1_nl;
  wire LOOPJ1_mux1h_2_nl;
  wire[4:0] LOOPJ1_mux1h_6_nl;
  wire LOOPJ1_mux1h_1_nl;
  wire mux_85_nl;
  wire mux_84_nl;
  wire mux_82_nl;
  wire mux_81_nl;
  wire[5:0] LOOPJ2_j_or_nl;
  wire[5:0] LOOPJ2_j_and_nl;
  wire[5:0] LOOPJ2_j_mux1h_nl;
  wire and_57_nl;
  wire and_59_nl;
  wire and_60_nl;
  wire and_61_nl;
  wire and_63_nl;
  wire and_65_nl;
  wire and_67_nl;
  wire and_68_nl;
  wire and_71_nl;
  wire and_74_nl;
  wire and_75_nl;
  wire and_76_nl;
  wire and_79_nl;
  wire and_81_nl;
  wire and_82_nl;
  wire and_83_nl;
  wire and_86_nl;
  wire and_88_nl;
  wire and_89_nl;
  wire and_90_nl;
  wire and_93_nl;
  wire and_95_nl;
  wire and_96_nl;
  wire and_97_nl;
  wire and_98_nl;
  wire and_99_nl;
  wire and_100_nl;
  wire and_101_nl;
  wire and_104_nl;
  wire and_107_nl;
  wire and_108_nl;
  wire and_109_nl;
  wire and_111_nl;
  wire and_113_nl;
  wire and_114_nl;
  wire and_115_nl;
  wire and_117_nl;
  wire and_119_nl;
  wire and_120_nl;
  wire and_121_nl;
  wire and_123_nl;
  wire and_125_nl;
  wire and_126_nl;
  wire and_127_nl;
  wire and_129_nl;
  wire and_131_nl;
  wire and_132_nl;
  wire and_133_nl;
  wire and_135_nl;
  wire and_137_nl;
  wire and_138_nl;
  wire and_139_nl;
  wire and_141_nl;
  wire and_143_nl;
  wire and_144_nl;
  wire and_145_nl;
  wire and_147_nl;
  wire and_149_nl;
  wire and_150_nl;
  wire and_151_nl;
  wire mux_89_nl;
  wire mux_88_nl;
  wire and_245_nl;
  wire mux_87_nl;
  wire mux_86_nl;
  wire or_463_nl;
  wire or_464_nl;
  wire or_465_nl;
  wire nor_58_nl;
  wire[5:0] LOOPJ2_j_or_1_nl;
  wire[5:0] LOOPJ2_j_and_1_nl;
  wire[5:0] LOOPJ2_j_mux1h_1_nl;
  wire LOOPJ1_nor_1_nl;
  wire mux_115_nl;
  wire mux_114_nl;
  wire mux_113_nl;
  wire mux_112_nl;
  wire mux_111_nl;
  wire or_318_nl;
  wire and_220_nl;
  wire mux_156_nl;
  wire mux_157_nl;
  wire nor_68_nl;
  wire and_288_nl;
  wire nor_69_nl;
  wire[1:0] LOOPI1_LOOPI1_and_1_nl;
  wire[1:0] LOOPI1_mux_1_nl;
  wire not_457_nl;
  wire[3:0] LOOPI1_mux1h_2_nl;
  wire and_301_nl;
  wire operator_7_false_operator_7_false_and_2_nl;
  wire operator_7_false_operator_7_false_and_3_nl;
  wire operator_7_false_mux_1_nl;
  wire operator_7_false_and_1_nl;
  wire operator_7_false_mux1h_4_nl;
  wire[3:0] operator_7_false_mux1h_5_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [1023:0] nl_ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_inst_q_chan1_rsci_idat;
  assign nl_ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_inst_q_chan1_rsci_idat
      = {q_chan1_rsci_idat_1023_1008 , q_chan1_rsci_idat_1007_992 , q_chan1_rsci_idat_991_976
      , q_chan1_rsci_idat_975_960 , q_chan1_rsci_idat_959_944 , q_chan1_rsci_idat_943_928
      , q_chan1_rsci_idat_927_912 , q_chan1_rsci_idat_911_896 , q_chan1_rsci_idat_895_880
      , q_chan1_rsci_idat_879_864 , q_chan1_rsci_idat_863_848 , q_chan1_rsci_idat_847_832
      , q_chan1_rsci_idat_831_816 , q_chan1_rsci_idat_815_800 , q_chan1_rsci_idat_799_784
      , q_chan1_rsci_idat_783_768 , q_chan1_rsci_idat_767_752 , q_chan1_rsci_idat_751_736
      , q_chan1_rsci_idat_735_720 , q_chan1_rsci_idat_719_704 , q_chan1_rsci_idat_703_688
      , q_chan1_rsci_idat_687_672 , q_chan1_rsci_idat_671_656 , q_chan1_rsci_idat_655_640
      , q_chan1_rsci_idat_639_624 , q_chan1_rsci_idat_623_608 , q_chan1_rsci_idat_607_592
      , q_chan1_rsci_idat_591_576 , q_chan1_rsci_idat_575_560 , q_chan1_rsci_idat_559_544
      , q_chan1_rsci_idat_543_528 , q_chan1_rsci_idat_527_512 , q_chan1_rsci_idat_511_496
      , q_chan1_rsci_idat_495_480 , q_chan1_rsci_idat_479_464 , q_chan1_rsci_idat_463_448
      , q_chan1_rsci_idat_447_432 , q_chan1_rsci_idat_431_416 , q_chan1_rsci_idat_415_400
      , q_chan1_rsci_idat_399_384 , q_chan1_rsci_idat_383_368 , q_chan1_rsci_idat_367_352
      , q_chan1_rsci_idat_351_336 , q_chan1_rsci_idat_335_320 , q_chan1_rsci_idat_319_304
      , q_chan1_rsci_idat_303_288 , q_chan1_rsci_idat_287_272 , q_chan1_rsci_idat_271_256
      , q_chan1_rsci_idat_255_240 , q_chan1_rsci_idat_239_224 , q_chan1_rsci_idat_223_208
      , q_chan1_rsci_idat_207_192 , q_chan1_rsci_idat_191_176 , q_chan1_rsci_idat_175_160
      , q_chan1_rsci_idat_159_144 , q_chan1_rsci_idat_143_128 , q_chan1_rsci_idat_127_112
      , q_chan1_rsci_idat_111_96 , q_chan1_rsci_idat_95_80 , q_chan1_rsci_idat_79_64
      , q_chan1_rsci_idat_63_48 , q_chan1_rsci_idat_47_32 , q_chan1_rsci_idat_31_16
      , q_chan1_rsci_idat_15_0};
  wire [1023:0] nl_ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_inst_k_chan1_rsci_idat;
  assign nl_ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_inst_k_chan1_rsci_idat
      = {k_chan1_rsci_idat_1023_1008 , k_chan1_rsci_idat_1007_992 , k_chan1_rsci_idat_991_976
      , k_chan1_rsci_idat_975_960 , k_chan1_rsci_idat_959_944 , k_chan1_rsci_idat_943_928
      , k_chan1_rsci_idat_927_912 , k_chan1_rsci_idat_911_896 , k_chan1_rsci_idat_895_880
      , k_chan1_rsci_idat_879_864 , k_chan1_rsci_idat_863_848 , k_chan1_rsci_idat_847_832
      , k_chan1_rsci_idat_831_816 , k_chan1_rsci_idat_815_800 , k_chan1_rsci_idat_799_784
      , k_chan1_rsci_idat_783_768 , k_chan1_rsci_idat_767_752 , k_chan1_rsci_idat_751_736
      , k_chan1_rsci_idat_735_720 , k_chan1_rsci_idat_719_704 , k_chan1_rsci_idat_703_688
      , k_chan1_rsci_idat_687_672 , k_chan1_rsci_idat_671_656 , k_chan1_rsci_idat_655_640
      , k_chan1_rsci_idat_639_624 , k_chan1_rsci_idat_623_608 , k_chan1_rsci_idat_607_592
      , k_chan1_rsci_idat_591_576 , k_chan1_rsci_idat_575_560 , k_chan1_rsci_idat_559_544
      , k_chan1_rsci_idat_543_528 , k_chan1_rsci_idat_527_512 , k_chan1_rsci_idat_511_496
      , k_chan1_rsci_idat_495_480 , k_chan1_rsci_idat_479_464 , k_chan1_rsci_idat_463_448
      , k_chan1_rsci_idat_447_432 , k_chan1_rsci_idat_431_416 , k_chan1_rsci_idat_415_400
      , k_chan1_rsci_idat_399_384 , k_chan1_rsci_idat_383_368 , k_chan1_rsci_idat_367_352
      , k_chan1_rsci_idat_351_336 , k_chan1_rsci_idat_335_320 , k_chan1_rsci_idat_319_304
      , k_chan1_rsci_idat_303_288 , k_chan1_rsci_idat_287_272 , k_chan1_rsci_idat_271_256
      , k_chan1_rsci_idat_255_240 , k_chan1_rsci_idat_239_224 , k_chan1_rsci_idat_223_208
      , k_chan1_rsci_idat_207_192 , k_chan1_rsci_idat_191_176 , k_chan1_rsci_idat_175_160
      , k_chan1_rsci_idat_159_144 , k_chan1_rsci_idat_143_128 , k_chan1_rsci_idat_127_112
      , k_chan1_rsci_idat_111_96 , k_chan1_rsci_idat_95_80 , k_chan1_rsci_idat_79_64
      , k_chan1_rsci_idat_63_48 , k_chan1_rsci_idat_47_32 , k_chan1_rsci_idat_31_16
      , k_chan1_rsci_idat_15_0};
  wire [1023:0] nl_ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_inst_v_chan1_rsci_idat;
  assign nl_ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_inst_v_chan1_rsci_idat
      = {v_chan1_rsci_idat_1023_1008 , v_chan1_rsci_idat_1007_992 , v_chan1_rsci_idat_991_976
      , v_chan1_rsci_idat_975_960 , v_chan1_rsci_idat_959_944 , v_chan1_rsci_idat_943_928
      , v_chan1_rsci_idat_927_912 , v_chan1_rsci_idat_911_896 , v_chan1_rsci_idat_895_880
      , v_chan1_rsci_idat_879_864 , v_chan1_rsci_idat_863_848 , v_chan1_rsci_idat_847_832
      , v_chan1_rsci_idat_831_816 , v_chan1_rsci_idat_815_800 , v_chan1_rsci_idat_799_784
      , v_chan1_rsci_idat_783_768 , v_chan1_rsci_idat_767_752 , v_chan1_rsci_idat_751_736
      , v_chan1_rsci_idat_735_720 , v_chan1_rsci_idat_719_704 , v_chan1_rsci_idat_703_688
      , v_chan1_rsci_idat_687_672 , v_chan1_rsci_idat_671_656 , v_chan1_rsci_idat_655_640
      , v_chan1_rsci_idat_639_624 , v_chan1_rsci_idat_623_608 , v_chan1_rsci_idat_607_592
      , v_chan1_rsci_idat_591_576 , v_chan1_rsci_idat_575_560 , v_chan1_rsci_idat_559_544
      , v_chan1_rsci_idat_543_528 , v_chan1_rsci_idat_527_512 , v_chan1_rsci_idat_511_496
      , v_chan1_rsci_idat_495_480 , v_chan1_rsci_idat_479_464 , v_chan1_rsci_idat_463_448
      , v_chan1_rsci_idat_447_432 , v_chan1_rsci_idat_431_416 , v_chan1_rsci_idat_415_400
      , v_chan1_rsci_idat_399_384 , v_chan1_rsci_idat_383_368 , v_chan1_rsci_idat_367_352
      , v_chan1_rsci_idat_351_336 , v_chan1_rsci_idat_335_320 , v_chan1_rsci_idat_319_304
      , v_chan1_rsci_idat_303_288 , v_chan1_rsci_idat_287_272 , v_chan1_rsci_idat_271_256
      , v_chan1_rsci_idat_255_240 , v_chan1_rsci_idat_239_224 , v_chan1_rsci_idat_223_208
      , v_chan1_rsci_idat_207_192 , v_chan1_rsci_idat_191_176 , v_chan1_rsci_idat_175_160
      , v_chan1_rsci_idat_159_144 , v_chan1_rsci_idat_143_128 , v_chan1_rsci_idat_127_112
      , v_chan1_rsci_idat_111_96 , v_chan1_rsci_idat_95_80 , v_chan1_rsci_idat_79_64
      , v_chan1_rsci_idat_63_48 , v_chan1_rsci_idat_47_32 , v_chan1_rsci_idat_31_16
      , v_chan1_rsci_idat_15_0};
  wire  nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_iswt0_pff;
  assign nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_iswt0_pff
      = ((or_111_cse | (fsm_output[3]) | or_145_cse) ^ (fsm_output[6])) & (fsm_output[8:7]==2'b00);
  wire  nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_oswt_1_pff;
  assign nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_oswt_1_pff
      = ~ mux_69_itm;
  wire  nl_ATTENTION_IP_Attention_Buffer_run_run_fsm_inst_LOOPJ2_C_66_tr0;
  assign nl_ATTENTION_IP_Attention_Buffer_run_run_fsm_inst_LOOPJ2_C_66_tr0 = ~((LOOPJ1_j_sva_5_0
      != (z_out_1[5:0])) | (z_out_1[6]));
  ATTENTION_IP_Attention_Buffer_run_din_chan_rsci ATTENTION_IP_Attention_Buffer_run_din_chan_rsci_inst
      (
      .din_chan_rsc_dat(din_chan_rsc_dat),
      .din_chan_rsc_vld(din_chan_rsc_vld),
      .din_chan_rsc_rdy(din_chan_rsc_rdy),
      .run_wen(run_wen),
      .din_chan_rsci_oswt(reg_din_chan_rsci_oswt_cse),
      .din_chan_rsci_wen_comp(din_chan_rsci_wen_comp),
      .din_chan_rsci_idat_mxwt(din_chan_rsci_idat_mxwt)
    );
  ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_inst
      (
      .q_chan1_rsc_dat(q_chan1_rsc_dat),
      .q_chan1_rsc_vld(q_chan1_rsc_vld),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy),
      .q_chan1_rsci_oswt(reg_q_chan1_rsci_oswt_cse),
      .q_chan1_rsci_wen_comp(q_chan1_rsci_wen_comp),
      .q_chan1_rsci_idat(nl_ATTENTION_IP_Attention_Buffer_run_q_chan1_rsci_inst_q_chan1_rsci_idat[1023:0])
    );
  ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_inst
      (
      .k_chan1_rsc_dat(k_chan1_rsc_dat),
      .k_chan1_rsc_vld(k_chan1_rsc_vld),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy),
      .k_chan1_rsci_oswt(reg_k_chan1_rsci_oswt_cse),
      .k_chan1_rsci_wen_comp(k_chan1_rsci_wen_comp),
      .k_chan1_rsci_idat(nl_ATTENTION_IP_Attention_Buffer_run_k_chan1_rsci_inst_k_chan1_rsci_idat[1023:0])
    );
  ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_inst
      (
      .v_chan1_rsc_dat(v_chan1_rsc_dat),
      .v_chan1_rsc_vld(v_chan1_rsc_vld),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy),
      .v_chan1_rsci_oswt(reg_v_chan1_rsci_oswt_cse),
      .v_chan1_rsci_wen_comp(v_chan1_rsci_wen_comp),
      .v_chan1_rsci_idat(nl_ATTENTION_IP_Attention_Buffer_run_v_chan1_rsci_inst_v_chan1_rsci_idat[1023:0])
    );
  ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1 ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .pp_buf_data_rsci_q_d(pp_buf_data_rsci_q_d),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .pp_buf_data_rsci_oswt_1(reg_pp_buf_data_rsci_oswt_1_cse),
      .pp_buf_data_rsci_q_d_mxwt(pp_buf_data_rsci_q_d_mxwt),
      .pp_buf_data_rsci_we_d_pff(pp_buf_data_rsci_we_d_iff),
      .pp_buf_data_rsci_iswt0_pff(nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_iswt0_pff),
      .pp_buf_data_rsci_re_d_pff(pp_buf_data_rsci_re_d_iff),
      .pp_buf_data_rsci_oswt_1_pff(nl_ATTENTION_IP_Attention_Buffer_run_pp_buf_data_rsci_1_inst_pp_buf_data_rsci_oswt_1_pff)
    );
  ATTENTION_IP_Attention_Buffer_run_staller ATTENTION_IP_Attention_Buffer_run_staller_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .run_wten(run_wten),
      .din_chan_rsci_wen_comp(din_chan_rsci_wen_comp),
      .q_chan1_rsci_wen_comp(q_chan1_rsci_wen_comp),
      .k_chan1_rsci_wen_comp(k_chan1_rsci_wen_comp),
      .v_chan1_rsci_wen_comp(v_chan1_rsci_wen_comp)
    );
  ATTENTION_IP_Attention_Buffer_run_run_fsm ATTENTION_IP_Attention_Buffer_run_run_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .LOOPK1_C_0_tr0(LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp),
      .LOOPJ1_C_64_tr0(LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp),
      .LOOPK2_C_65_tr0(LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm),
      .LOOPK3_C_65_tr0(LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm),
      .LOOPJ2_C_66_tr0(nl_ATTENTION_IP_Attention_Buffer_run_run_fsm_inst_LOOPJ2_C_66_tr0),
      .LOOPI1_C_0_tr0(LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp)
    );
  assign LOOPK3_and_cse = run_wen & (~(or_dcpl_104 | (fsm_output[2:1]!=2'b11) | or_dcpl_101));
  assign LOOPK2_and_cse = run_wen & (~(or_dcpl_109 | (fsm_output[2:1]!=2'b10) | or_dcpl_101));
  assign LOOPJ2_and_cse = run_wen & (~(or_dcpl_114 | (fsm_output[2:1]!=2'b01) | or_dcpl_101));
  assign or_108_cse = (fsm_output[4:3]!=2'b00);
  assign or_146_cse_1 = (~ (fsm_output[6])) | (fsm_output[8]);
  assign or_145_cse = (fsm_output[5:4]!=2'b00);
  assign or_111_cse = (fsm_output[2:1]!=2'b00);
  assign nor_28_cse = ~((fsm_output[0]) | (fsm_output[5]));
  assign channel_in_data_and_cse = run_wen & (~(or_dcpl_113 | (fsm_output[7]) | or_111_cse
      | or_dcpl_101));
  assign mux_65_nl = MUX_s_1_2_2(mux_16_cse, mux_tmp_59, fsm_output[2]);
  assign mux_66_nl = MUX_s_1_2_2(mux_65_nl, mux_tmp_62, fsm_output[1]);
  assign mux_67_nl = MUX_s_1_2_2(mux_66_nl, or_tmp_23, or_108_cse);
  assign mux_60_nl = MUX_s_1_2_2(mux_tmp_59, or_tmp_23, fsm_output[2]);
  assign mux_63_nl = MUX_s_1_2_2(mux_tmp_62, mux_60_nl, fsm_output[1]);
  assign mux_64_nl = MUX_s_1_2_2(mux_63_nl, or_tmp_23, or_108_cse);
  assign mux_68_nl = MUX_s_1_2_2(mux_67_nl, mux_64_nl, fsm_output[0]);
  assign mux_69_itm = MUX_s_1_2_2(mux_68_nl, or_tmp_23, fsm_output[5]);
  assign and_237_cse = (fsm_output[2:1]==2'b11);
  assign nor_49_cse = ~((fsm_output[1:0]!=2'b00));
  assign nor_53_cse = ~(mux_tmp_102 | (fsm_output[0]));
  assign nor_54_cse = ~(mux_tmp_104 | (fsm_output[0]));
  assign or_319_cse = (fsm_output[4:1]!=4'b0000);
  assign or_158_cse_1 = (fsm_output[5:3]!=3'b000);
  assign or_478_cse = (~ (fsm_output[8])) | (fsm_output[6]);
  assign or_472_cse = (fsm_output[8:7]!=2'b01);
  assign or_476_cse = (~ (fsm_output[8])) | (fsm_output[1]) | (fsm_output[6]);
  assign nl_LOOPK1_acc_1_tmp = LOOPJ1_acc_itm_6_0 + 7'b0000001;
  assign LOOPK1_acc_1_tmp = nl_LOOPK1_acc_1_tmp[6:0];
  assign nl_LOOPK2_acc_tmp_sva_mx0w2 = conv_u2u_6_7(length) + conv_u2u_6_7(LOOPK2_acc_1_itm);
  assign LOOPK2_acc_tmp_sva_mx0w2 = nl_LOOPK2_acc_tmp_sva_mx0w2[6:0];
  assign nl_LOOPK3_acc_psp_sva_mx0w4 = conv_u2u_6_7(length) + conv_u2u_5_7(LOOPK2_acc_1_itm[5:1]);
  assign LOOPK3_acc_psp_sva_mx0w4 = nl_LOOPK3_acc_psp_sva_mx0w4[6:0];
  assign nl_operator_6_false_acc_psp_sva_1 = conv_s2s_7_9({(z_out_1[5:0]) , (length[0])})
      + conv_u2s_7_9({length , 1'b1});
  assign operator_6_false_acc_psp_sva_1 = nl_operator_6_false_acc_psp_sva_1[8:0];
  assign LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp = ~((LOOPI1_i_sva != (z_out_1[3:0]))
      | (z_out_1[4]));
  assign LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp = ~((({LOOPJ1_j_sva_7 , LOOPJ1_j_sva_6
      , LOOPJ1_j_sva_5_0}) != (operator_6_false_acc_psp_sva_1[7:0])) | (operator_6_false_acc_psp_sva_1[8]));
  assign LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp = ~((LOOPJ1_acc_itm_6_0 != (z_out_1[6:0]))
      | (z_out_1[7]));
  assign or_dcpl = ~((LOOPK1_acc_1_tmp[2:1]==2'b11));
  assign or_dcpl_1 = or_dcpl | (~ (LOOPK1_acc_1_tmp[0]));
  assign or_dcpl_2 = ~((LOOPK1_acc_1_tmp[4:3]==2'b11));
  assign or_dcpl_3 = LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp | (~ (LOOPK1_acc_1_tmp[5]));
  assign or_dcpl_4 = or_dcpl_3 | or_dcpl_2;
  assign or_dcpl_6 = or_dcpl | (LOOPK1_acc_1_tmp[0]);
  assign or_dcpl_8 = (LOOPK1_acc_1_tmp[2:1]!=2'b00);
  assign or_dcpl_9 = or_dcpl_8 | (~ (LOOPK1_acc_1_tmp[0]));
  assign or_dcpl_10 = (LOOPK1_acc_1_tmp[4:3]!=2'b00);
  assign or_dcpl_11 = LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp | (LOOPK1_acc_1_tmp[5]);
  assign or_dcpl_12 = or_dcpl_11 | or_dcpl_10;
  assign or_dcpl_14 = (LOOPK1_acc_1_tmp[2:1]!=2'b10);
  assign or_dcpl_15 = or_dcpl_14 | (~ (LOOPK1_acc_1_tmp[0]));
  assign or_dcpl_17 = (LOOPK1_acc_1_tmp[2:1]!=2'b01);
  assign or_dcpl_18 = or_dcpl_17 | (LOOPK1_acc_1_tmp[0]);
  assign or_dcpl_20 = or_dcpl_14 | (LOOPK1_acc_1_tmp[0]);
  assign or_dcpl_22 = or_dcpl_17 | (~ (LOOPK1_acc_1_tmp[0]));
  assign or_dcpl_30 = or_dcpl_8 | (LOOPK1_acc_1_tmp[0]);
  assign or_dcpl_33 = (LOOPK1_acc_1_tmp[4:3]!=2'b10);
  assign or_dcpl_34 = or_dcpl_3 | or_dcpl_33;
  assign or_dcpl_36 = (LOOPK1_acc_1_tmp[4:3]!=2'b01);
  assign or_dcpl_37 = or_dcpl_11 | or_dcpl_36;
  assign or_dcpl_53 = or_dcpl_3 | or_dcpl_36;
  assign or_dcpl_55 = or_dcpl_11 | or_dcpl_33;
  assign or_dcpl_71 = or_dcpl_3 | or_dcpl_10;
  assign or_dcpl_73 = or_dcpl_11 | or_dcpl_2;
  assign mux_16_cse = MUX_s_1_2_2(or_478_cse, (fsm_output[8]), fsm_output[7]);
  assign and_dcpl_7 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_8 = and_dcpl_7 & nor_28_cse;
  assign and_dcpl_9 = ~((fsm_output[2:1]!=2'b00));
  assign and_dcpl_10 = ~((fsm_output[8]) | (fsm_output[6]));
  assign and_dcpl_11 = and_dcpl_10 & (~ (fsm_output[7]));
  assign and_dcpl_12 = and_dcpl_11 & and_dcpl_9;
  assign and_dcpl_14 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_15 = and_dcpl_14 & nor_28_cse;
  assign and_dcpl_16 = (fsm_output[2:1]==2'b01);
  assign and_dcpl_18 = (fsm_output[8:6]==3'b100);
  assign or_dcpl_93 = (fsm_output[0]) | (fsm_output[5]);
  assign or_dcpl_99 = (~ (fsm_output[0])) | (fsm_output[5]);
  assign or_dcpl_101 = or_108_cse | or_dcpl_99;
  assign or_dcpl_104 = or_478_cse | (fsm_output[7]);
  assign or_dcpl_109 = or_146_cse_1 | (~ (fsm_output[7]));
  assign or_dcpl_113 = (fsm_output[8]) | (fsm_output[6]);
  assign or_dcpl_114 = or_dcpl_113 | (~ (fsm_output[7]));
  assign and_dcpl_23 = (~ (fsm_output[8])) & (fsm_output[6]);
  assign and_dcpl_24 = and_dcpl_23 & (~ (fsm_output[7]));
  assign nor_34_cse = ~((fsm_output[7:6]!=2'b00));
  assign or_tmp_23 = nor_34_cse | (fsm_output[8]);
  assign or_143_nl = (fsm_output[7:6]!=2'b00);
  assign mux_tmp_26 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), or_143_nl);
  assign mux_tmp_27 = MUX_s_1_2_2(mux_tmp_26, or_tmp_23, or_111_cse);
  assign mux_29_nl = MUX_s_1_2_2(mux_16_cse, mux_tmp_26, or_111_cse);
  assign mux_30_nl = MUX_s_1_2_2(mux_29_nl, mux_tmp_27, fsm_output[3]);
  assign mux_tmp_31 = MUX_s_1_2_2(mux_30_nl, or_tmp_23, fsm_output[4]);
  assign mux_32_nl = MUX_s_1_2_2(mux_16_cse, mux_tmp_26, fsm_output[2]);
  assign mux_33_nl = MUX_s_1_2_2(mux_32_nl, mux_tmp_27, fsm_output[3]);
  assign mux_tmp_34 = MUX_s_1_2_2(mux_33_nl, or_tmp_23, fsm_output[4]);
  assign and_dcpl_32 = (fsm_output[0]) & (~ (fsm_output[5]));
  assign and_dcpl_33 = and_dcpl_7 & and_dcpl_32;
  assign and_dcpl_34 = and_dcpl_12 & and_dcpl_33;
  assign and_dcpl_35 = (fsm_output[2:1]==2'b10);
  assign and_dcpl_36 = and_dcpl_10 & (fsm_output[7]);
  assign and_dcpl_38 = and_dcpl_36 & and_dcpl_35 & and_dcpl_33;
  assign and_dcpl_40 = and_dcpl_23 & (fsm_output[7]);
  assign and_dcpl_42 = and_dcpl_40 & and_237_cse & and_dcpl_33;
  assign or_dcpl_121 = ~((LOOPJ1_acc_itm_6_0[3]) & (LOOPJ1_acc_itm_6_0[5]));
  assign or_dcpl_122 = or_dcpl_121 | (~ (LOOPJ1_acc_itm_6_0[4]));
  assign or_dcpl_123 = ~((LOOPJ1_acc_itm_6_0[1:0]==2'b11));
  assign or_dcpl_124 = or_dcpl_123 | (~ (LOOPJ1_acc_itm_6_0[2]));
  assign or_dcpl_126 = (LOOPJ1_acc_itm_6_0[1:0]!=2'b10);
  assign or_dcpl_127 = or_dcpl_126 | (~ (LOOPJ1_acc_itm_6_0[2]));
  assign or_dcpl_129 = (LOOPJ1_acc_itm_6_0[3]) | (LOOPJ1_acc_itm_6_0[5]);
  assign or_dcpl_130 = or_dcpl_129 | (LOOPJ1_acc_itm_6_0[4]);
  assign or_dcpl_131 = (LOOPJ1_acc_itm_6_0[1:0]!=2'b01);
  assign or_dcpl_132 = or_dcpl_131 | (LOOPJ1_acc_itm_6_0[2]);
  assign or_dcpl_134 = or_dcpl_131 | (~ (LOOPJ1_acc_itm_6_0[2]));
  assign or_dcpl_136 = or_dcpl_126 | (LOOPJ1_acc_itm_6_0[2]);
  assign or_dcpl_138 = (LOOPJ1_acc_itm_6_0[1:0]!=2'b00);
  assign or_dcpl_139 = or_dcpl_138 | (~ (LOOPJ1_acc_itm_6_0[2]));
  assign or_dcpl_141 = or_dcpl_123 | (LOOPJ1_acc_itm_6_0[2]);
  assign or_dcpl_149 = or_dcpl_138 | (LOOPJ1_acc_itm_6_0[2]);
  assign or_dcpl_152 = (LOOPJ1_acc_itm_6_0[3]) | (~ (LOOPJ1_acc_itm_6_0[5]));
  assign or_dcpl_153 = or_dcpl_152 | (~ (LOOPJ1_acc_itm_6_0[4]));
  assign or_dcpl_155 = (~ (LOOPJ1_acc_itm_6_0[3])) | (LOOPJ1_acc_itm_6_0[5]);
  assign or_dcpl_156 = or_dcpl_155 | (LOOPJ1_acc_itm_6_0[4]);
  assign or_dcpl_172 = or_dcpl_121 | (LOOPJ1_acc_itm_6_0[4]);
  assign or_dcpl_174 = or_dcpl_129 | (~ (LOOPJ1_acc_itm_6_0[4]));
  assign or_dcpl_190 = or_dcpl_152 | (LOOPJ1_acc_itm_6_0[4]);
  assign or_dcpl_192 = or_dcpl_155 | (~ (LOOPJ1_acc_itm_6_0[4]));
  assign or_tmp_46 = (~ (fsm_output[1])) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_tmp_53 = MUX_s_1_2_2(or_dcpl_113, or_146_cse_1, fsm_output[1]);
  assign mux_tmp_58 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[6]);
  assign mux_tmp_59 = MUX_s_1_2_2(mux_tmp_58, or_146_cse_1, fsm_output[7]);
  assign mux_61_nl = MUX_s_1_2_2(mux_tmp_58, or_dcpl_113, fsm_output[7]);
  assign mux_tmp_62 = MUX_s_1_2_2(mux_16_cse, mux_61_nl, fsm_output[2]);
  assign or_tmp_51 = (fsm_output[7:6]!=2'b01);
  assign or_tmp_53 = (fsm_output[7:6]!=2'b10);
  assign or_268_nl = (fsm_output[4:2]!=3'b000);
  assign mux_71_nl = MUX_s_1_2_2(or_tmp_53, or_tmp_51, or_268_nl);
  assign mux_70_nl = MUX_s_1_2_2(or_tmp_53, or_tmp_51, or_319_cse);
  assign mux_72_nl = MUX_s_1_2_2(mux_71_nl, mux_70_nl, fsm_output[0]);
  assign mux_73_nl = MUX_s_1_2_2(mux_72_nl, or_tmp_51, fsm_output[5]);
  assign and_dcpl_51 = ~(mux_73_nl | (fsm_output[8]));
  assign mux_tmp_74 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[2]);
  assign mux_77_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), and_237_cse);
  assign mux_78_nl = MUX_s_1_2_2(mux_77_nl, (fsm_output[6]), or_108_cse);
  assign or_270_nl = (fsm_output[2]) | (~ (fsm_output[6]));
  assign mux_75_nl = MUX_s_1_2_2(or_270_nl, mux_tmp_74, fsm_output[1]);
  assign mux_76_nl = MUX_s_1_2_2(mux_75_nl, (fsm_output[6]), or_108_cse);
  assign mux_79_nl = MUX_s_1_2_2(mux_78_nl, mux_76_nl, fsm_output[0]);
  assign mux_80_nl = MUX_s_1_2_2(mux_79_nl, (fsm_output[6]), fsm_output[5]);
  assign and_dcpl_53 = (~ mux_80_nl) & (fsm_output[8:7]==2'b01);
  assign mux_tmp_83 = MUX_s_1_2_2(or_dcpl_104, or_dcpl_109, or_108_cse);
  assign and_dcpl_54 = ~((fsm_output[8]) | (fsm_output[4]));
  assign and_dcpl_55 = and_dcpl_54 & nor_28_cse;
  assign nor_tmp_13 = (fsm_output[7:6]==2'b11);
  assign or_tmp_70 = (~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign or_286_nl = (~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[6]));
  assign mux_tmp_90 = MUX_s_1_2_2(or_286_nl, or_tmp_70, fsm_output[1]);
  assign or_283_nl = (fsm_output[2:1]!=2'b00) | (~ nor_tmp_13);
  assign mux_tmp_91 = MUX_s_1_2_2(mux_tmp_90, or_283_nl, fsm_output[3]);
  assign and_dcpl_57 = and_dcpl_54 & and_dcpl_32;
  assign or_tmp_74 = (fsm_output[2]) | (~ (fsm_output[7])) | (fsm_output[6]);
  assign or_287_nl = (fsm_output[2]) | (~ nor_tmp_13);
  assign mux_tmp_92 = MUX_s_1_2_2(or_tmp_74, or_287_nl, fsm_output[1]);
  assign nand_12_nl = ~((fsm_output[1]) & (fsm_output[2]) & (~ (fsm_output[7])) &
      (fsm_output[6]));
  assign mux_tmp_93 = MUX_s_1_2_2(nand_12_nl, mux_tmp_92, fsm_output[3]);
  assign mux_tmp_94 = MUX_s_1_2_2((~ or_tmp_51), nor_tmp_13, fsm_output[2]);
  assign mux_tmp_95 = MUX_s_1_2_2((~ mux_tmp_94), or_tmp_74, fsm_output[1]);
  assign and_dcpl_61 = ~(mux_tmp_95 | (fsm_output[8]));
  assign and_dcpl_63 = and_dcpl_14 & and_dcpl_32;
  assign mux_tmp_96 = MUX_s_1_2_2((~ or_tmp_70), mux_tmp_94, fsm_output[1]);
  assign and_dcpl_65 = mux_tmp_96 & (~ (fsm_output[8]));
  assign and_dcpl_68 = ~((fsm_output[8]) | (fsm_output[0]));
  assign and_dcpl_69 = and_dcpl_68 & (~ (fsm_output[5]));
  assign nand_nl = ~((fsm_output[3]) & (~ mux_tmp_90));
  assign or_292_nl = (fsm_output[3:1]!=3'b000) | (~ nor_tmp_13);
  assign mux_tmp_97 = MUX_s_1_2_2(nand_nl, or_292_nl, fsm_output[4]);
  assign and_dcpl_71 = (~ (fsm_output[8])) & (fsm_output[0]);
  assign and_dcpl_72 = and_dcpl_71 & (~ (fsm_output[5]));
  assign nand_14_nl = ~((fsm_output[3]) & (fsm_output[1]) & (fsm_output[2]) & (~
      (fsm_output[7])) & (fsm_output[6]));
  assign or_293_nl = (fsm_output[3]) | mux_tmp_92;
  assign mux_tmp_98 = MUX_s_1_2_2(nand_14_nl, or_293_nl, fsm_output[4]);
  assign and_dcpl_76 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_77 = and_dcpl_76 & nor_28_cse;
  assign and_dcpl_79 = and_dcpl_76 & and_dcpl_32;
  assign and_dcpl_83 = (~ (fsm_output[8])) & (fsm_output[4]);
  assign and_dcpl_84 = and_dcpl_83 & nor_28_cse;
  assign and_dcpl_86 = and_dcpl_83 & and_dcpl_32;
  assign and_dcpl_90 = (fsm_output[4:3]==2'b11);
  assign and_dcpl_91 = and_dcpl_90 & nor_28_cse;
  assign and_dcpl_93 = and_dcpl_90 & and_dcpl_32;
  assign nand_1_nl = ~((fsm_output[4:3]==2'b11) & (~ mux_tmp_90));
  assign or_297_nl = (fsm_output[4:1]!=4'b0000) | (~ nor_tmp_13);
  assign mux_tmp_99 = MUX_s_1_2_2(nand_1_nl, or_297_nl, fsm_output[5]);
  assign nand_16_nl = ~((fsm_output[4]) & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[2])
      & (~ (fsm_output[7])) & (fsm_output[6]));
  assign or_299_nl = (fsm_output[4:3]!=2'b00) | mux_tmp_92;
  assign mux_tmp_100 = MUX_s_1_2_2(nand_16_nl, or_299_nl, fsm_output[5]);
  assign and_dcpl_101 = (~ (fsm_output[0])) & (fsm_output[5]);
  assign and_dcpl_102 = and_dcpl_7 & and_dcpl_101;
  assign and_dcpl_104 = (fsm_output[0]) & (fsm_output[5]);
  assign and_dcpl_105 = and_dcpl_7 & and_dcpl_104;
  assign and_dcpl_109 = and_dcpl_54 & and_dcpl_101;
  assign and_dcpl_111 = and_dcpl_54 & and_dcpl_104;
  assign and_dcpl_115 = and_dcpl_14 & and_dcpl_101;
  assign and_dcpl_117 = and_dcpl_14 & and_dcpl_104;
  assign and_dcpl_121 = and_dcpl_68 & (fsm_output[5]);
  assign and_dcpl_123 = and_dcpl_71 & (fsm_output[5]);
  assign and_dcpl_127 = and_dcpl_76 & and_dcpl_101;
  assign and_dcpl_129 = and_dcpl_76 & and_dcpl_104;
  assign and_dcpl_133 = and_dcpl_83 & and_dcpl_101;
  assign and_dcpl_135 = and_dcpl_83 & and_dcpl_104;
  assign and_dcpl_139 = and_dcpl_90 & and_dcpl_101;
  assign and_dcpl_141 = and_dcpl_90 & and_dcpl_104;
  assign or_305_nl = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[1]) | (fsm_output[2])
      | (fsm_output[7]) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign nor_40_nl = ~((~ (fsm_output[2])) | (fsm_output[7]) | (~ (fsm_output[6]))
      | (fsm_output[8]));
  assign nor_41_nl = ~((~ (fsm_output[2])) | (~ (fsm_output[7])) | (fsm_output[6])
      | (fsm_output[8]));
  assign mux_101_nl = MUX_s_1_2_2(nor_40_nl, nor_41_nl, fsm_output[1]);
  assign nand_2_nl = ~((fsm_output[4:3]==2'b11) & mux_101_nl);
  assign mux_tmp_102 = MUX_s_1_2_2(or_305_nl, nand_2_nl, fsm_output[5]);
  assign or_tmp_96 = (fsm_output[2]) | (~ (fsm_output[7])) | (~ (fsm_output[6]))
      | (fsm_output[8]);
  assign or_309_nl = (fsm_output[2]) | (fsm_output[7]) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_103_nl = MUX_s_1_2_2(or_tmp_96, or_309_nl, fsm_output[1]);
  assign or_311_nl = (fsm_output[4:3]!=2'b00) | mux_103_nl;
  assign nand_17_nl = ~((fsm_output[4]) & (fsm_output[3]) & (fsm_output[1]) & (fsm_output[2])
      & (~ (fsm_output[7])) & (fsm_output[6]) & (~ (fsm_output[8])));
  assign mux_tmp_104 = MUX_s_1_2_2(or_311_nl, nand_17_nl, fsm_output[5]);
  assign mux_tmp_105 = MUX_s_1_2_2(or_dcpl_114, or_dcpl_104, fsm_output[2]);
  assign mux_tmp_106 = MUX_s_1_2_2(mux_tmp_105, or_tmp_96, fsm_output[1]);
  assign nand_18_nl = ~((fsm_output[2]) & (fsm_output[7]) & (fsm_output[6]) & (~
      (fsm_output[8])));
  assign mux_107_nl = MUX_s_1_2_2(nand_18_nl, mux_tmp_105, fsm_output[1]);
  assign and_dcpl_151 = (~ mux_107_nl) & and_dcpl_8;
  assign and_dcpl_152 = and_dcpl_11 & and_dcpl_16;
  assign and_dcpl_153 = and_dcpl_152 & and_dcpl_8;
  assign and_dcpl_154 = and_dcpl_11 & and_dcpl_35;
  assign and_dcpl_155 = and_dcpl_154 & and_dcpl_8;
  assign and_dcpl_156 = and_dcpl_154 & and_dcpl_33;
  assign and_dcpl_157 = and_dcpl_11 & and_237_cse;
  assign and_dcpl_158 = and_dcpl_157 & and_dcpl_8;
  assign and_dcpl_159 = and_dcpl_157 & and_dcpl_33;
  assign and_dcpl_160 = and_dcpl_12 & and_dcpl_15;
  assign and_dcpl_161 = and_dcpl_12 & and_dcpl_63;
  assign and_dcpl_162 = and_dcpl_152 & and_dcpl_15;
  assign and_dcpl_163 = and_dcpl_152 & and_dcpl_63;
  assign and_dcpl_164 = and_dcpl_154 & and_dcpl_15;
  assign and_dcpl_165 = and_dcpl_154 & and_dcpl_63;
  assign and_dcpl_166 = and_dcpl_157 & and_dcpl_15;
  assign and_dcpl_167 = and_dcpl_157 & and_dcpl_63;
  assign and_dcpl_168 = and_dcpl_12 & and_dcpl_77;
  assign and_dcpl_169 = and_dcpl_12 & and_dcpl_79;
  assign and_dcpl_170 = and_dcpl_152 & and_dcpl_77;
  assign and_dcpl_171 = and_dcpl_152 & and_dcpl_79;
  assign and_dcpl_172 = and_dcpl_154 & and_dcpl_77;
  assign and_dcpl_173 = and_dcpl_154 & and_dcpl_79;
  assign and_dcpl_174 = and_dcpl_157 & and_dcpl_77;
  assign and_dcpl_175 = and_dcpl_157 & and_dcpl_79;
  assign and_dcpl_176 = and_dcpl_12 & and_dcpl_91;
  assign and_dcpl_177 = and_dcpl_12 & and_dcpl_93;
  assign and_dcpl_178 = and_dcpl_152 & and_dcpl_91;
  assign and_dcpl_179 = and_dcpl_152 & and_dcpl_93;
  assign and_dcpl_180 = and_dcpl_154 & and_dcpl_91;
  assign and_dcpl_181 = and_dcpl_154 & and_dcpl_93;
  assign and_dcpl_182 = and_dcpl_157 & and_dcpl_91;
  assign and_dcpl_183 = and_dcpl_157 & and_dcpl_93;
  assign and_dcpl_184 = and_dcpl_12 & and_dcpl_102;
  assign and_dcpl_185 = and_dcpl_12 & and_dcpl_105;
  assign and_dcpl_186 = and_dcpl_152 & and_dcpl_102;
  assign and_dcpl_187 = and_dcpl_152 & and_dcpl_105;
  assign and_dcpl_188 = and_dcpl_154 & and_dcpl_102;
  assign and_dcpl_189 = and_dcpl_154 & and_dcpl_105;
  assign and_dcpl_190 = and_dcpl_157 & and_dcpl_102;
  assign and_dcpl_191 = and_dcpl_157 & and_dcpl_105;
  assign and_dcpl_192 = and_dcpl_12 & and_dcpl_115;
  assign and_dcpl_193 = and_dcpl_12 & and_dcpl_117;
  assign and_dcpl_194 = and_dcpl_152 & and_dcpl_115;
  assign and_dcpl_195 = and_dcpl_152 & and_dcpl_117;
  assign and_dcpl_196 = and_dcpl_154 & and_dcpl_115;
  assign and_dcpl_197 = and_dcpl_154 & and_dcpl_117;
  assign and_dcpl_198 = and_dcpl_157 & and_dcpl_115;
  assign and_dcpl_199 = and_dcpl_157 & and_dcpl_117;
  assign and_dcpl_200 = and_dcpl_12 & and_dcpl_127;
  assign and_dcpl_201 = and_dcpl_12 & and_dcpl_129;
  assign and_dcpl_202 = and_dcpl_152 & and_dcpl_127;
  assign and_dcpl_203 = and_dcpl_152 & and_dcpl_129;
  assign and_dcpl_204 = and_dcpl_154 & and_dcpl_127;
  assign and_dcpl_205 = and_dcpl_154 & and_dcpl_129;
  assign and_dcpl_206 = and_dcpl_157 & and_dcpl_127;
  assign and_dcpl_207 = and_dcpl_157 & and_dcpl_129;
  assign and_dcpl_208 = and_dcpl_12 & and_dcpl_139;
  assign and_dcpl_209 = and_dcpl_12 & and_dcpl_141;
  assign and_dcpl_210 = and_dcpl_152 & and_dcpl_139;
  assign and_dcpl_211 = and_dcpl_152 & and_dcpl_141;
  assign and_dcpl_212 = and_dcpl_154 & and_dcpl_139;
  assign and_dcpl_213 = and_dcpl_154 & and_dcpl_141;
  assign and_dcpl_214 = and_dcpl_157 & and_dcpl_139;
  assign and_dcpl_215 = and_dcpl_157 & and_dcpl_141;
  assign and_dcpl_216 = and_dcpl_24 & and_dcpl_9;
  assign and_dcpl_217 = and_dcpl_216 & and_dcpl_8;
  assign and_dcpl_218 = and_dcpl_216 & and_dcpl_33;
  assign or_dcpl_219 = (fsm_output[8]) | (fsm_output[4]);
  assign or_dcpl_220 = or_dcpl_219 | or_dcpl_93;
  assign or_dcpl_222 = or_dcpl_219 | or_dcpl_99;
  assign or_dcpl_226 = (fsm_output[4:3]!=2'b01);
  assign or_dcpl_227 = or_dcpl_226 | or_dcpl_93;
  assign or_dcpl_228 = mux_tmp_95 | (fsm_output[8]);
  assign or_dcpl_230 = or_dcpl_226 | or_dcpl_99;
  assign or_dcpl_232 = (~ mux_tmp_96) | (fsm_output[8]);
  assign or_dcpl_235 = (fsm_output[8]) | (fsm_output[0]);
  assign or_dcpl_236 = or_dcpl_235 | (fsm_output[5]);
  assign or_dcpl_238 = (fsm_output[8]) | (~ (fsm_output[0]));
  assign or_dcpl_239 = or_dcpl_238 | (fsm_output[5]);
  assign or_dcpl_243 = (fsm_output[4:3]!=2'b10);
  assign or_dcpl_244 = or_dcpl_243 | or_dcpl_93;
  assign or_dcpl_246 = or_dcpl_243 | or_dcpl_99;
  assign or_dcpl_250 = (fsm_output[8]) | (~ (fsm_output[4]));
  assign or_dcpl_251 = or_dcpl_250 | or_dcpl_93;
  assign or_dcpl_253 = or_dcpl_250 | or_dcpl_99;
  assign or_dcpl_257 = ~((fsm_output[4:3]==2'b11));
  assign or_dcpl_258 = or_dcpl_257 | or_dcpl_93;
  assign or_dcpl_260 = or_dcpl_257 | or_dcpl_99;
  assign or_dcpl_268 = (fsm_output[0]) | (~ (fsm_output[5]));
  assign or_dcpl_269 = or_108_cse | or_dcpl_268;
  assign or_dcpl_271 = ~((fsm_output[0]) & (fsm_output[5]));
  assign or_dcpl_272 = or_108_cse | or_dcpl_271;
  assign or_dcpl_276 = or_dcpl_219 | or_dcpl_268;
  assign or_dcpl_278 = or_dcpl_219 | or_dcpl_271;
  assign or_dcpl_282 = or_dcpl_226 | or_dcpl_268;
  assign or_dcpl_284 = or_dcpl_226 | or_dcpl_271;
  assign or_dcpl_288 = or_dcpl_235 | (~ (fsm_output[5]));
  assign or_dcpl_290 = or_dcpl_238 | (~ (fsm_output[5]));
  assign or_dcpl_294 = or_dcpl_243 | or_dcpl_268;
  assign or_dcpl_296 = or_dcpl_243 | or_dcpl_271;
  assign or_dcpl_300 = or_dcpl_250 | or_dcpl_268;
  assign or_dcpl_302 = or_dcpl_250 | or_dcpl_271;
  assign or_dcpl_306 = or_dcpl_257 | or_dcpl_268;
  assign or_dcpl_308 = or_dcpl_257 | or_dcpl_271;
  assign mux_tmp_140 = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[7]);
  assign or_453_nl = (fsm_output[8:7]!=2'b10);
  assign mux_tmp_143 = MUX_s_1_2_2(or_453_nl, or_472_cse, fsm_output[6]);
  assign LOOPI1_i_sva_mx0c0 = and_dcpl_12 & and_dcpl_8;
  assign or_141_nl = (fsm_output[0]) | LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp;
  assign mux_35_nl = MUX_s_1_2_2(mux_tmp_34, mux_tmp_31, or_141_nl);
  assign mux_36_itm = MUX_s_1_2_2(mux_35_nl, or_tmp_23, fsm_output[5]);
  assign nor_33_nl = ~((fsm_output[1]) | (fsm_output[8]));
  assign and_nl = (fsm_output[1]) & (fsm_output[8]);
  assign mux_25_nl = MUX_s_1_2_2(nor_33_nl, and_nl, fsm_output[3]);
  assign LOOPJ1_j_sva_mx0c2 = mux_25_nl & nor_34_cse & (~((fsm_output[2]) | (fsm_output[4])))
      & nor_28_cse;
  assign or_105_nl = and_237_cse | (fsm_output[8:6]!=3'b100);
  assign mux_108_nl = MUX_s_1_2_2(or_105_nl, or_dcpl_109, or_108_cse);
  assign mux_109_nl = MUX_s_1_2_2(mux_tmp_83, mux_108_nl, fsm_output[0]);
  assign mux_110_itm = MUX_s_1_2_2(mux_109_nl, or_dcpl_109, fsm_output[5]);
  assign LOOPJ1_j_and_ssc = run_wen & ((and_dcpl_24 & and_dcpl_16 & and_dcpl_7 &
      (~ LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp) & nor_28_cse) | (~ mux_36_itm) | LOOPJ1_j_sva_mx0c2);
  assign nl_LOOPJ1_acc_sdt = ({LOOPJ1_j_sva_7 , LOOPJ1_j_sva_6 , LOOPJ1_j_sva_5_0})
      + 8'b00000001;
  assign LOOPJ1_acc_sdt = nl_LOOPJ1_acc_sdt[7:0];
  assign nor_145_cse = ~((fsm_output[5:4]!=2'b00));
  assign LOOPJ1_mux_nl = MUX_s_1_2_2((LOOPJ1_acc_itm_6_0[6]), (LOOPK3_acc_psp_sva_mx0w4[6]),
      mux_110_itm);
  assign LOOPJ1_LOOPJ1_and_nl = LOOPJ1_mux_nl & (~(and_dcpl_51 | and_dcpl_38 | and_dcpl_53));
  assign LOOPJ1_mux1h_2_nl = MUX1HOT_s_1_4_2((LOOPK2_acc_tmp_sva_mx0w2[6]), (LOOPJ1_acc_itm_6_0[6]),
      (LOOPK3_acc_psp_sva_mx0w4[5]), (LOOPJ1_acc_itm_6_0[5]), {and_dcpl_38 , and_dcpl_53
      , and_dcpl_42 , (~ mux_110_itm)});
  assign LOOPJ1_and_1_nl = LOOPJ1_mux1h_2_nl & (~ and_dcpl_51);
  assign LOOPJ1_mux1h_6_nl = MUX1HOT_v_5_5_2((LOOPJ1_j_sva_5_0[5:1]), (LOOPK2_acc_tmp_sva_mx0w2[5:1]),
      (LOOPJ1_acc_itm_6_0[5:1]), (LOOPK3_acc_psp_sva_mx0w4[4:0]), (LOOPJ1_acc_itm_6_0[4:0]),
      {and_dcpl_51 , and_dcpl_38 , and_dcpl_53 , and_dcpl_42 , (~ mux_110_itm)});
  assign mux_81_nl = MUX_s_1_2_2(or_dcpl_104, or_dcpl_109, and_237_cse);
  assign mux_82_nl = MUX_s_1_2_2(mux_81_nl, or_dcpl_109, or_108_cse);
  assign mux_84_nl = MUX_s_1_2_2(mux_tmp_83, mux_82_nl, fsm_output[0]);
  assign mux_85_nl = MUX_s_1_2_2(mux_84_nl, or_dcpl_109, fsm_output[5]);
  assign LOOPJ1_mux1h_1_nl = MUX1HOT_s_1_4_2((LOOPJ1_j_sva_5_0[0]), (LOOPK2_acc_tmp_sva_mx0w2[0]),
      (LOOPJ1_acc_itm_6_0[0]), (LOOPK2_acc_1_itm[0]), {and_dcpl_51 , and_dcpl_38
      , and_dcpl_53 , (~ mux_85_nl)});
  assign and_57_nl = (~ mux_tmp_91) & and_dcpl_55;
  assign and_59_nl = (~ mux_tmp_91) & and_dcpl_57;
  assign and_60_nl = (~ mux_tmp_93) & and_dcpl_55;
  assign and_61_nl = (~ mux_tmp_93) & and_dcpl_57;
  assign and_63_nl = and_dcpl_61 & and_dcpl_15;
  assign and_65_nl = and_dcpl_61 & and_dcpl_63;
  assign and_67_nl = and_dcpl_65 & and_dcpl_15;
  assign and_68_nl = and_dcpl_65 & and_dcpl_63;
  assign and_71_nl = (~ mux_tmp_97) & and_dcpl_69;
  assign and_74_nl = (~ mux_tmp_97) & and_dcpl_72;
  assign and_75_nl = (~ mux_tmp_98) & and_dcpl_69;
  assign and_76_nl = (~ mux_tmp_98) & and_dcpl_72;
  assign and_79_nl = and_dcpl_61 & and_dcpl_77;
  assign and_81_nl = and_dcpl_61 & and_dcpl_79;
  assign and_82_nl = and_dcpl_65 & and_dcpl_77;
  assign and_83_nl = and_dcpl_65 & and_dcpl_79;
  assign and_86_nl = (~ mux_tmp_91) & and_dcpl_84;
  assign and_88_nl = (~ mux_tmp_91) & and_dcpl_86;
  assign and_89_nl = (~ mux_tmp_93) & and_dcpl_84;
  assign and_90_nl = (~ mux_tmp_93) & and_dcpl_86;
  assign and_93_nl = and_dcpl_61 & and_dcpl_91;
  assign and_95_nl = and_dcpl_61 & and_dcpl_93;
  assign and_96_nl = and_dcpl_65 & and_dcpl_91;
  assign and_97_nl = and_dcpl_65 & and_dcpl_93;
  assign and_98_nl = (~ mux_tmp_99) & and_dcpl_68;
  assign and_99_nl = (~ mux_tmp_99) & and_dcpl_71;
  assign and_100_nl = (~ mux_tmp_100) & and_dcpl_68;
  assign and_101_nl = (~ mux_tmp_100) & and_dcpl_71;
  assign and_104_nl = and_dcpl_61 & and_dcpl_102;
  assign and_107_nl = and_dcpl_61 & and_dcpl_105;
  assign and_108_nl = and_dcpl_65 & and_dcpl_102;
  assign and_109_nl = and_dcpl_65 & and_dcpl_105;
  assign and_111_nl = (~ mux_tmp_91) & and_dcpl_109;
  assign and_113_nl = (~ mux_tmp_91) & and_dcpl_111;
  assign and_114_nl = (~ mux_tmp_93) & and_dcpl_109;
  assign and_115_nl = (~ mux_tmp_93) & and_dcpl_111;
  assign and_117_nl = and_dcpl_61 & and_dcpl_115;
  assign and_119_nl = and_dcpl_61 & and_dcpl_117;
  assign and_120_nl = and_dcpl_65 & and_dcpl_115;
  assign and_121_nl = and_dcpl_65 & and_dcpl_117;
  assign and_123_nl = (~ mux_tmp_97) & and_dcpl_121;
  assign and_125_nl = (~ mux_tmp_97) & and_dcpl_123;
  assign and_126_nl = (~ mux_tmp_98) & and_dcpl_121;
  assign and_127_nl = (~ mux_tmp_98) & and_dcpl_123;
  assign and_129_nl = and_dcpl_61 & and_dcpl_127;
  assign and_131_nl = and_dcpl_61 & and_dcpl_129;
  assign and_132_nl = and_dcpl_65 & and_dcpl_127;
  assign and_133_nl = and_dcpl_65 & and_dcpl_129;
  assign and_135_nl = (~ mux_tmp_91) & and_dcpl_133;
  assign and_137_nl = (~ mux_tmp_91) & and_dcpl_135;
  assign and_138_nl = (~ mux_tmp_93) & and_dcpl_133;
  assign and_139_nl = (~ mux_tmp_93) & and_dcpl_135;
  assign and_141_nl = and_dcpl_61 & and_dcpl_139;
  assign and_143_nl = and_dcpl_61 & and_dcpl_141;
  assign and_144_nl = and_dcpl_65 & and_dcpl_139;
  assign and_145_nl = and_dcpl_65 & and_dcpl_141;
  assign and_147_nl = (~ mux_tmp_102) & (fsm_output[0]);
  assign and_149_nl = (~ mux_tmp_104) & (fsm_output[0]);
  assign and_150_nl = (~ mux_tmp_106) & and_dcpl_8;
  assign and_151_nl = (~ mux_tmp_106) & and_dcpl_33;
  assign LOOPJ2_j_mux1h_nl = MUX1HOT_v_6_62_2(6'b000001, 6'b000010, 6'b000011, 6'b000100,
      6'b000101, 6'b000110, 6'b000111, 6'b001000, 6'b001001, 6'b001010, 6'b001011,
      6'b001100, 6'b001101, 6'b001110, 6'b001111, 6'b010000, 6'b010001, 6'b010010,
      6'b010011, 6'b010100, 6'b010101, 6'b010110, 6'b010111, 6'b011000, 6'b011001,
      6'b011010, 6'b011011, 6'b011100, 6'b011101, 6'b011110, 6'b011111, 6'b100000,
      6'b100001, 6'b100010, 6'b100011, 6'b100100, 6'b100101, 6'b100110, 6'b100111,
      6'b101000, 6'b101001, 6'b101010, 6'b101011, 6'b101100, 6'b101101, 6'b101110,
      6'b101111, 6'b110000, 6'b110001, 6'b110010, 6'b110011, 6'b110100, 6'b110101,
      6'b110110, 6'b110111, 6'b111000, 6'b111001, 6'b111010, 6'b111011, 6'b111100,
      6'b111101, 6'b111110, {and_57_nl , and_59_nl , and_60_nl , and_61_nl , and_63_nl
      , and_65_nl , and_67_nl , and_68_nl , and_71_nl , and_74_nl , and_75_nl , and_76_nl
      , and_79_nl , and_81_nl , and_82_nl , and_83_nl , and_86_nl , and_88_nl , and_89_nl
      , and_90_nl , and_93_nl , and_95_nl , and_96_nl , and_97_nl , and_98_nl , and_99_nl
      , and_100_nl , and_101_nl , and_104_nl , and_107_nl , and_108_nl , and_109_nl
      , and_111_nl , and_113_nl , and_114_nl , and_115_nl , and_117_nl , and_119_nl
      , and_120_nl , and_121_nl , and_123_nl , and_125_nl , and_126_nl , and_127_nl
      , and_129_nl , and_131_nl , and_132_nl , and_133_nl , and_135_nl , and_137_nl
      , and_138_nl , and_139_nl , and_141_nl , and_143_nl , and_144_nl , and_145_nl
      , nor_53_cse , and_147_nl , nor_54_cse , and_149_nl , and_150_nl , and_151_nl});
  assign and_245_nl = (fsm_output[6]) & ((fsm_output[5:2]!=4'b0000));
  assign or_463_nl = (fsm_output[5:2]!=4'b0001);
  assign or_464_nl = (~ (fsm_output[0])) | (fsm_output[2]) | (fsm_output[3]) | (fsm_output[4])
      | (fsm_output[5]);
  assign mux_86_nl = MUX_s_1_2_2(or_463_nl, or_464_nl, fsm_output[1]);
  assign or_465_nl = nor_49_cse | (fsm_output[5:2]!=4'b0001);
  assign mux_87_nl = MUX_s_1_2_2(mux_86_nl, or_465_nl, fsm_output[6]);
  assign mux_88_nl = MUX_s_1_2_2(and_245_nl, mux_87_nl, fsm_output[7]);
  assign nor_58_nl = ~((fsm_output[7:6]!=2'b00) | ((fsm_output[2:0]==3'b111)) | (fsm_output[5:3]!=3'b000));
  assign mux_89_nl = MUX_s_1_2_2(mux_88_nl, nor_58_nl, fsm_output[8]);
  assign LOOPJ2_j_and_nl = MUX_v_6_2_2(6'b000000, LOOPJ2_j_mux1h_nl, mux_89_nl);
  assign LOOPJ2_j_or_nl = MUX_v_6_2_2(LOOPJ2_j_and_nl, 6'b111111, and_dcpl_151);
  assign pp_buf_data_rsci_radr_d = {LOOPJ1_LOOPJ1_and_nl , LOOPJ1_and_1_nl , LOOPJ1_mux1h_6_nl
      , LOOPJ1_mux1h_1_nl , LOOPJ2_j_or_nl};
  assign LOOPJ2_j_mux1h_1_nl = MUX1HOT_v_6_62_2(6'b111110, 6'b000001, 6'b111101,
      6'b000010, 6'b111100, 6'b000011, 6'b111011, 6'b000100, 6'b111010, 6'b000101,
      6'b111001, 6'b000110, 6'b111000, 6'b000111, 6'b110111, 6'b001000, 6'b110110,
      6'b001001, 6'b110101, 6'b001010, 6'b110100, 6'b001011, 6'b110011, 6'b001100,
      6'b110010, 6'b001101, 6'b110001, 6'b001110, 6'b110000, 6'b001111, 6'b101111,
      6'b010000, 6'b101110, 6'b010001, 6'b101101, 6'b010010, 6'b101100, 6'b010011,
      6'b101011, 6'b010100, 6'b101010, 6'b010101, 6'b101001, 6'b010110, 6'b101000,
      6'b010111, 6'b100111, 6'b011000, 6'b100110, 6'b011001, 6'b100101, 6'b011010,
      6'b100100, 6'b011011, 6'b100011, 6'b011100, 6'b100010, 6'b011101, 6'b100001,
      6'b011110, 6'b100000, 6'b011111, {and_dcpl_155 , and_dcpl_156 , and_dcpl_158
      , and_dcpl_159 , and_dcpl_160 , and_dcpl_161 , and_dcpl_162 , and_dcpl_163
      , and_dcpl_164 , and_dcpl_165 , and_dcpl_166 , and_dcpl_167 , and_dcpl_168
      , and_dcpl_169 , and_dcpl_170 , and_dcpl_171 , and_dcpl_172 , and_dcpl_173
      , and_dcpl_174 , and_dcpl_175 , and_dcpl_176 , and_dcpl_177 , and_dcpl_178
      , and_dcpl_179 , and_dcpl_180 , and_dcpl_181 , and_dcpl_182 , and_dcpl_183
      , and_dcpl_184 , and_dcpl_185 , and_dcpl_186 , and_dcpl_187 , and_dcpl_188
      , and_dcpl_189 , and_dcpl_190 , and_dcpl_191 , and_dcpl_192 , and_dcpl_193
      , and_dcpl_194 , and_dcpl_195 , and_dcpl_196 , and_dcpl_197 , and_dcpl_198
      , and_dcpl_199 , and_dcpl_200 , and_dcpl_201 , and_dcpl_202 , and_dcpl_203
      , and_dcpl_204 , and_dcpl_205 , and_dcpl_206 , and_dcpl_207 , and_dcpl_208
      , and_dcpl_209 , and_dcpl_210 , and_dcpl_211 , and_dcpl_212 , and_dcpl_213
      , and_dcpl_214 , and_dcpl_215 , and_dcpl_217 , and_dcpl_218});
  assign mux_113_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), or_319_cse);
  assign or_318_nl = (~ (fsm_output[2])) | (fsm_output[6]);
  assign mux_111_nl = MUX_s_1_2_2(mux_tmp_74, or_318_nl, fsm_output[1]);
  assign mux_112_nl = MUX_s_1_2_2(mux_111_nl, (fsm_output[6]), or_108_cse);
  assign mux_114_nl = MUX_s_1_2_2(mux_113_nl, mux_112_nl, fsm_output[0]);
  assign mux_115_nl = MUX_s_1_2_2(mux_114_nl, (fsm_output[6]), fsm_output[5]);
  assign LOOPJ1_nor_1_nl = ~(mux_115_nl | (fsm_output[8:7]!=2'b00));
  assign LOOPJ2_j_and_1_nl = MUX_v_6_2_2(6'b000000, LOOPJ2_j_mux1h_1_nl, LOOPJ1_nor_1_nl);
  assign LOOPJ2_j_or_1_nl = MUX_v_6_2_2(LOOPJ2_j_and_1_nl, 6'b111111, and_dcpl_153);
  assign pp_buf_data_rsci_wadr_d = {LOOPJ1_j_sva_7 , LOOPJ1_j_sva_6 , LOOPJ1_j_sva_5_0
      , LOOPJ2_j_or_1_nl};
  assign and_220_nl = and_dcpl_152 & and_dcpl_33;
  assign pp_buf_data_rsci_d_d = MUX1HOT_v_16_64_2(channel_in_data_63_lpi_4, LOOPJ2_asn_itm,
      channel_in_data_62_lpi_4, channel_in_data_1_lpi_4, channel_in_data_61_lpi_4,
      channel_in_data_2_lpi_4, channel_in_data_60_lpi_4, channel_in_data_3_lpi_4,
      channel_in_data_59_lpi_4, channel_in_data_4_lpi_4, channel_in_data_58_lpi_4,
      channel_in_data_5_lpi_4, channel_in_data_57_lpi_4, channel_in_data_6_lpi_4,
      channel_in_data_56_lpi_4, channel_in_data_7_lpi_4, channel_in_data_55_lpi_4,
      channel_in_data_8_lpi_4, channel_in_data_54_lpi_4, channel_in_data_9_lpi_4,
      channel_in_data_53_lpi_4, channel_in_data_10_lpi_4, channel_in_data_52_lpi_4,
      channel_in_data_11_lpi_4, channel_in_data_51_lpi_4, channel_in_data_12_lpi_4,
      channel_in_data_50_lpi_4, channel_in_data_13_lpi_4, channel_in_data_49_lpi_4,
      channel_in_data_14_lpi_4, channel_in_data_48_lpi_4, channel_in_data_15_lpi_4,
      channel_in_data_47_lpi_4, channel_in_data_16_lpi_4, channel_in_data_46_lpi_4,
      channel_in_data_17_lpi_4, channel_in_data_45_lpi_4, channel_in_data_18_lpi_4,
      channel_in_data_44_lpi_4, channel_in_data_19_lpi_4, channel_in_data_43_lpi_4,
      channel_in_data_20_lpi_4, channel_in_data_42_lpi_4, channel_in_data_21_lpi_4,
      channel_in_data_41_lpi_4, channel_in_data_22_lpi_4, channel_in_data_40_lpi_4,
      channel_in_data_23_lpi_4, channel_in_data_39_lpi_4, channel_in_data_24_lpi_4,
      channel_in_data_38_lpi_4, channel_in_data_25_lpi_4, channel_in_data_37_lpi_4,
      channel_in_data_26_lpi_4, channel_in_data_36_lpi_4, channel_in_data_27_lpi_4,
      channel_in_data_35_lpi_4, channel_in_data_28_lpi_4, channel_in_data_34_lpi_4,
      channel_in_data_29_lpi_4, channel_in_data_33_lpi_4, channel_in_data_30_lpi_4,
      channel_in_data_32_lpi_4, channel_in_data_31_lpi_4, {and_dcpl_153 , and_220_nl
      , and_dcpl_155 , and_dcpl_156 , and_dcpl_158 , and_dcpl_159 , and_dcpl_160
      , and_dcpl_161 , and_dcpl_162 , and_dcpl_163 , and_dcpl_164 , and_dcpl_165
      , and_dcpl_166 , and_dcpl_167 , and_dcpl_168 , and_dcpl_169 , and_dcpl_170
      , and_dcpl_171 , and_dcpl_172 , and_dcpl_173 , and_dcpl_174 , and_dcpl_175
      , and_dcpl_176 , and_dcpl_177 , and_dcpl_178 , and_dcpl_179 , and_dcpl_180
      , and_dcpl_181 , and_dcpl_182 , and_dcpl_183 , and_dcpl_184 , and_dcpl_185
      , and_dcpl_186 , and_dcpl_187 , and_dcpl_188 , and_dcpl_189 , and_dcpl_190
      , and_dcpl_191 , and_dcpl_192 , and_dcpl_193 , and_dcpl_194 , and_dcpl_195
      , and_dcpl_196 , and_dcpl_197 , and_dcpl_198 , and_dcpl_199 , and_dcpl_200
      , and_dcpl_201 , and_dcpl_202 , and_dcpl_203 , and_dcpl_204 , and_dcpl_205
      , and_dcpl_206 , and_dcpl_207 , and_dcpl_208 , and_dcpl_209 , and_dcpl_210
      , and_dcpl_211 , and_dcpl_212 , and_dcpl_213 , and_dcpl_214 , and_dcpl_215
      , and_dcpl_217 , and_dcpl_218});
  assign pp_buf_data_rsci_we_d_pff = pp_buf_data_rsci_we_d_iff;
  assign pp_buf_data_rsci_re_d_pff = pp_buf_data_rsci_re_d_iff;
  assign and_dcpl = (~ (fsm_output[6])) & (fsm_output[8]);
  assign and_dcpl_227 = nor_145_cse & (fsm_output[3]);
  assign and_dcpl_246 = ~((fsm_output[5:3]!=3'b000));
  assign nor_63_cse = ~((fsm_output[0]) | (fsm_output[7]));
  assign and_252_itm = and_dcpl_227 & (fsm_output[2:1]==2'b01) & nor_63_cse & and_dcpl;
  assign and_263_itm = and_dcpl_227 & and_dcpl_9 & (fsm_output[0]) & (~ (fsm_output[7]))
      & and_dcpl;
  assign and_271_itm = and_dcpl_246 & and_dcpl_9 & (fsm_output[0]) & (~ (fsm_output[7]))
      & and_dcpl_10;
  assign and_277_itm = and_dcpl_246 & and_dcpl_16 & nor_63_cse & (fsm_output[6])
      & (~ (fsm_output[8]));
  assign nor_68_nl = ~((~ (fsm_output[7])) | (fsm_output[1]) | (~ (fsm_output[2]))
      | (fsm_output[3]));
  assign and_288_nl = (fsm_output[7]) & (fsm_output[1]) & (fsm_output[2]) & (~ (fsm_output[3]));
  assign mux_157_nl = MUX_s_1_2_2(nor_68_nl, and_288_nl, fsm_output[6]);
  assign nor_69_nl = ~((fsm_output[6]) | (fsm_output[7]) | (fsm_output[1]) | (fsm_output[2])
      | (~ (fsm_output[3])));
  assign mux_156_nl = MUX_s_1_2_2(mux_157_nl, nor_69_nl, fsm_output[8]);
  assign and_280_itm = mux_156_nl & nor_145_cse & (fsm_output[0]);
  assign and_286_itm = (fsm_output[5:3]==3'b001) & and_dcpl_16 & nor_63_cse & (~
      (fsm_output[6])) & (fsm_output[8]);
  always @(posedge clk) begin
    if ( run_wen & (LOOPI1_i_sva_mx0c0 | (and_dcpl_18 & and_dcpl_16 & and_dcpl_15))
        ) begin
      LOOPI1_i_sva <= MUX_v_4_2_2(4'b0000, (z_out[3:0]), LOOPI1_i_not_1_nl);
    end
  end
  always @(posedge clk) begin
    if ( LOOPK3_and_cse ) begin
      v_chan1_rsci_idat_511_496 <= LOOPJ2_asn_itm_31;
      v_chan1_rsci_idat_527_512 <= LOOPJ2_asn_itm_30;
      v_chan1_rsci_idat_495_480 <= LOOPJ2_asn_itm_32;
      v_chan1_rsci_idat_543_528 <= LOOPJ2_asn_itm_29;
      v_chan1_rsci_idat_479_464 <= LOOPJ2_asn_itm_33;
      v_chan1_rsci_idat_559_544 <= LOOPJ2_asn_itm_28;
      v_chan1_rsci_idat_463_448 <= LOOPJ2_asn_itm_34;
      v_chan1_rsci_idat_575_560 <= LOOPJ2_asn_itm_27;
      v_chan1_rsci_idat_447_432 <= LOOPJ2_asn_itm_35;
      v_chan1_rsci_idat_591_576 <= LOOPJ2_asn_itm_26;
      v_chan1_rsci_idat_431_416 <= LOOPJ2_asn_itm_36;
      v_chan1_rsci_idat_607_592 <= LOOPJ2_asn_itm_25;
      v_chan1_rsci_idat_415_400 <= LOOPJ2_asn_itm_37;
      v_chan1_rsci_idat_623_608 <= LOOPJ2_asn_itm_24;
      v_chan1_rsci_idat_399_384 <= LOOPJ2_asn_itm_38;
      v_chan1_rsci_idat_639_624 <= LOOPJ2_asn_itm_23;
      v_chan1_rsci_idat_383_368 <= LOOPJ2_asn_itm_39;
      v_chan1_rsci_idat_655_640 <= LOOPJ2_asn_itm_22;
      v_chan1_rsci_idat_367_352 <= LOOPJ2_asn_itm_40;
      v_chan1_rsci_idat_671_656 <= LOOPJ2_asn_itm_21;
      v_chan1_rsci_idat_351_336 <= LOOPJ2_asn_itm_41;
      v_chan1_rsci_idat_687_672 <= LOOPJ2_asn_itm_20;
      v_chan1_rsci_idat_335_320 <= LOOPJ2_asn_itm_42;
      v_chan1_rsci_idat_703_688 <= LOOPJ2_asn_itm_19;
      v_chan1_rsci_idat_319_304 <= LOOPJ2_asn_itm_43;
      v_chan1_rsci_idat_719_704 <= LOOPJ2_asn_itm_18;
      v_chan1_rsci_idat_303_288 <= LOOPJ2_asn_itm_44;
      v_chan1_rsci_idat_735_720 <= LOOPJ2_asn_itm_17;
      v_chan1_rsci_idat_287_272 <= LOOPJ2_asn_itm_45;
      v_chan1_rsci_idat_751_736 <= LOOPJ2_asn_itm_16;
      v_chan1_rsci_idat_271_256 <= LOOPJ2_asn_itm_46;
      v_chan1_rsci_idat_767_752 <= LOOPJ2_asn_itm_15;
      v_chan1_rsci_idat_255_240 <= LOOPJ2_asn_itm_47;
      v_chan1_rsci_idat_783_768 <= LOOPJ2_asn_itm_14;
      v_chan1_rsci_idat_239_224 <= LOOPJ2_asn_itm_48;
      v_chan1_rsci_idat_799_784 <= LOOPJ2_asn_itm_13;
      v_chan1_rsci_idat_223_208 <= LOOPJ2_asn_itm_49;
      v_chan1_rsci_idat_815_800 <= LOOPJ2_asn_itm_12;
      v_chan1_rsci_idat_207_192 <= LOOPJ2_asn_itm_50;
      v_chan1_rsci_idat_831_816 <= LOOPJ2_asn_itm_11;
      v_chan1_rsci_idat_191_176 <= LOOPJ2_asn_itm_51;
      v_chan1_rsci_idat_847_832 <= LOOPJ2_asn_itm_10;
      v_chan1_rsci_idat_175_160 <= LOOPJ2_asn_itm_52;
      v_chan1_rsci_idat_863_848 <= LOOPJ2_asn_itm_9;
      v_chan1_rsci_idat_159_144 <= LOOPJ2_asn_itm_53;
      v_chan1_rsci_idat_879_864 <= LOOPJ2_asn_itm_8;
      v_chan1_rsci_idat_143_128 <= LOOPJ2_asn_itm_54;
      v_chan1_rsci_idat_895_880 <= LOOPJ2_asn_itm_7;
      v_chan1_rsci_idat_127_112 <= LOOPJ2_asn_itm_55;
      v_chan1_rsci_idat_911_896 <= LOOPJ2_asn_itm_6;
      v_chan1_rsci_idat_111_96 <= LOOPJ2_asn_itm_56;
      v_chan1_rsci_idat_927_912 <= LOOPJ2_asn_itm_5;
      v_chan1_rsci_idat_95_80 <= LOOPJ2_asn_itm_57;
      v_chan1_rsci_idat_943_928 <= LOOPJ2_asn_itm_4;
      v_chan1_rsci_idat_79_64 <= LOOPJ2_asn_itm_58;
      v_chan1_rsci_idat_959_944 <= LOOPJ2_asn_itm_3;
      v_chan1_rsci_idat_63_48 <= LOOPJ2_asn_itm_59;
      v_chan1_rsci_idat_975_960 <= LOOPJ2_asn_itm_2;
      v_chan1_rsci_idat_47_32 <= LOOPJ2_asn_itm_60;
      v_chan1_rsci_idat_991_976 <= LOOPJ2_asn_itm_1;
      v_chan1_rsci_idat_31_16 <= LOOPJ2_asn_itm_61;
      v_chan1_rsci_idat_1007_992 <= LOOPJ2_asn_itm;
      v_chan1_rsci_idat_15_0 <= LOOPJ2_asn_itm_62;
      v_chan1_rsci_idat_1023_1008 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( LOOPK2_and_cse ) begin
      k_chan1_rsci_idat_511_496 <= LOOPJ2_asn_itm_31;
      k_chan1_rsci_idat_527_512 <= LOOPJ2_asn_itm_30;
      k_chan1_rsci_idat_495_480 <= LOOPJ2_asn_itm_32;
      k_chan1_rsci_idat_543_528 <= LOOPJ2_asn_itm_29;
      k_chan1_rsci_idat_479_464 <= LOOPJ2_asn_itm_33;
      k_chan1_rsci_idat_559_544 <= LOOPJ2_asn_itm_28;
      k_chan1_rsci_idat_463_448 <= LOOPJ2_asn_itm_34;
      k_chan1_rsci_idat_575_560 <= LOOPJ2_asn_itm_27;
      k_chan1_rsci_idat_447_432 <= LOOPJ2_asn_itm_35;
      k_chan1_rsci_idat_591_576 <= LOOPJ2_asn_itm_26;
      k_chan1_rsci_idat_431_416 <= LOOPJ2_asn_itm_36;
      k_chan1_rsci_idat_607_592 <= LOOPJ2_asn_itm_25;
      k_chan1_rsci_idat_415_400 <= LOOPJ2_asn_itm_37;
      k_chan1_rsci_idat_623_608 <= LOOPJ2_asn_itm_24;
      k_chan1_rsci_idat_399_384 <= LOOPJ2_asn_itm_38;
      k_chan1_rsci_idat_639_624 <= LOOPJ2_asn_itm_23;
      k_chan1_rsci_idat_383_368 <= LOOPJ2_asn_itm_39;
      k_chan1_rsci_idat_655_640 <= LOOPJ2_asn_itm_22;
      k_chan1_rsci_idat_367_352 <= LOOPJ2_asn_itm_40;
      k_chan1_rsci_idat_671_656 <= LOOPJ2_asn_itm_21;
      k_chan1_rsci_idat_351_336 <= LOOPJ2_asn_itm_41;
      k_chan1_rsci_idat_687_672 <= LOOPJ2_asn_itm_20;
      k_chan1_rsci_idat_335_320 <= LOOPJ2_asn_itm_42;
      k_chan1_rsci_idat_703_688 <= LOOPJ2_asn_itm_19;
      k_chan1_rsci_idat_319_304 <= LOOPJ2_asn_itm_43;
      k_chan1_rsci_idat_719_704 <= LOOPJ2_asn_itm_18;
      k_chan1_rsci_idat_303_288 <= LOOPJ2_asn_itm_44;
      k_chan1_rsci_idat_735_720 <= LOOPJ2_asn_itm_17;
      k_chan1_rsci_idat_287_272 <= LOOPJ2_asn_itm_45;
      k_chan1_rsci_idat_751_736 <= LOOPJ2_asn_itm_16;
      k_chan1_rsci_idat_271_256 <= LOOPJ2_asn_itm_46;
      k_chan1_rsci_idat_767_752 <= LOOPJ2_asn_itm_15;
      k_chan1_rsci_idat_255_240 <= LOOPJ2_asn_itm_47;
      k_chan1_rsci_idat_783_768 <= LOOPJ2_asn_itm_14;
      k_chan1_rsci_idat_239_224 <= LOOPJ2_asn_itm_48;
      k_chan1_rsci_idat_799_784 <= LOOPJ2_asn_itm_13;
      k_chan1_rsci_idat_223_208 <= LOOPJ2_asn_itm_49;
      k_chan1_rsci_idat_815_800 <= LOOPJ2_asn_itm_12;
      k_chan1_rsci_idat_207_192 <= LOOPJ2_asn_itm_50;
      k_chan1_rsci_idat_831_816 <= LOOPJ2_asn_itm_11;
      k_chan1_rsci_idat_191_176 <= LOOPJ2_asn_itm_51;
      k_chan1_rsci_idat_847_832 <= LOOPJ2_asn_itm_10;
      k_chan1_rsci_idat_175_160 <= LOOPJ2_asn_itm_52;
      k_chan1_rsci_idat_863_848 <= LOOPJ2_asn_itm_9;
      k_chan1_rsci_idat_159_144 <= LOOPJ2_asn_itm_53;
      k_chan1_rsci_idat_879_864 <= LOOPJ2_asn_itm_8;
      k_chan1_rsci_idat_143_128 <= LOOPJ2_asn_itm_54;
      k_chan1_rsci_idat_895_880 <= LOOPJ2_asn_itm_7;
      k_chan1_rsci_idat_127_112 <= LOOPJ2_asn_itm_55;
      k_chan1_rsci_idat_911_896 <= LOOPJ2_asn_itm_6;
      k_chan1_rsci_idat_111_96 <= LOOPJ2_asn_itm_56;
      k_chan1_rsci_idat_927_912 <= LOOPJ2_asn_itm_5;
      k_chan1_rsci_idat_95_80 <= LOOPJ2_asn_itm_57;
      k_chan1_rsci_idat_943_928 <= LOOPJ2_asn_itm_4;
      k_chan1_rsci_idat_79_64 <= LOOPJ2_asn_itm_58;
      k_chan1_rsci_idat_959_944 <= LOOPJ2_asn_itm_3;
      k_chan1_rsci_idat_63_48 <= LOOPJ2_asn_itm_59;
      k_chan1_rsci_idat_975_960 <= LOOPJ2_asn_itm_2;
      k_chan1_rsci_idat_47_32 <= LOOPJ2_asn_itm_60;
      k_chan1_rsci_idat_991_976 <= LOOPJ2_asn_itm_1;
      k_chan1_rsci_idat_31_16 <= LOOPJ2_asn_itm_61;
      k_chan1_rsci_idat_1007_992 <= LOOPJ2_asn_itm;
      k_chan1_rsci_idat_15_0 <= LOOPJ2_asn_itm_62;
      k_chan1_rsci_idat_1023_1008 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( LOOPJ2_and_cse ) begin
      q_chan1_rsci_idat_511_496 <= LOOPJ2_asn_itm_31;
      q_chan1_rsci_idat_527_512 <= LOOPJ2_asn_itm_30;
      q_chan1_rsci_idat_495_480 <= LOOPJ2_asn_itm_32;
      q_chan1_rsci_idat_543_528 <= LOOPJ2_asn_itm_29;
      q_chan1_rsci_idat_479_464 <= LOOPJ2_asn_itm_33;
      q_chan1_rsci_idat_559_544 <= LOOPJ2_asn_itm_28;
      q_chan1_rsci_idat_463_448 <= LOOPJ2_asn_itm_34;
      q_chan1_rsci_idat_575_560 <= LOOPJ2_asn_itm_27;
      q_chan1_rsci_idat_447_432 <= LOOPJ2_asn_itm_35;
      q_chan1_rsci_idat_591_576 <= LOOPJ2_asn_itm_26;
      q_chan1_rsci_idat_431_416 <= LOOPJ2_asn_itm_36;
      q_chan1_rsci_idat_607_592 <= LOOPJ2_asn_itm_25;
      q_chan1_rsci_idat_415_400 <= LOOPJ2_asn_itm_37;
      q_chan1_rsci_idat_623_608 <= LOOPJ2_asn_itm_24;
      q_chan1_rsci_idat_399_384 <= LOOPJ2_asn_itm_38;
      q_chan1_rsci_idat_639_624 <= LOOPJ2_asn_itm_23;
      q_chan1_rsci_idat_383_368 <= LOOPJ2_asn_itm_39;
      q_chan1_rsci_idat_655_640 <= LOOPJ2_asn_itm_22;
      q_chan1_rsci_idat_367_352 <= LOOPJ2_asn_itm_40;
      q_chan1_rsci_idat_671_656 <= LOOPJ2_asn_itm_21;
      q_chan1_rsci_idat_351_336 <= LOOPJ2_asn_itm_41;
      q_chan1_rsci_idat_687_672 <= LOOPJ2_asn_itm_20;
      q_chan1_rsci_idat_335_320 <= LOOPJ2_asn_itm_42;
      q_chan1_rsci_idat_703_688 <= LOOPJ2_asn_itm_19;
      q_chan1_rsci_idat_319_304 <= LOOPJ2_asn_itm_43;
      q_chan1_rsci_idat_719_704 <= LOOPJ2_asn_itm_18;
      q_chan1_rsci_idat_303_288 <= LOOPJ2_asn_itm_44;
      q_chan1_rsci_idat_735_720 <= LOOPJ2_asn_itm_17;
      q_chan1_rsci_idat_287_272 <= LOOPJ2_asn_itm_45;
      q_chan1_rsci_idat_751_736 <= LOOPJ2_asn_itm_16;
      q_chan1_rsci_idat_271_256 <= LOOPJ2_asn_itm_46;
      q_chan1_rsci_idat_767_752 <= LOOPJ2_asn_itm_15;
      q_chan1_rsci_idat_255_240 <= LOOPJ2_asn_itm_47;
      q_chan1_rsci_idat_783_768 <= LOOPJ2_asn_itm_14;
      q_chan1_rsci_idat_239_224 <= LOOPJ2_asn_itm_48;
      q_chan1_rsci_idat_799_784 <= LOOPJ2_asn_itm_13;
      q_chan1_rsci_idat_223_208 <= LOOPJ2_asn_itm_49;
      q_chan1_rsci_idat_815_800 <= LOOPJ2_asn_itm_12;
      q_chan1_rsci_idat_207_192 <= LOOPJ2_asn_itm_50;
      q_chan1_rsci_idat_831_816 <= LOOPJ2_asn_itm_11;
      q_chan1_rsci_idat_191_176 <= LOOPJ2_asn_itm_51;
      q_chan1_rsci_idat_847_832 <= LOOPJ2_asn_itm_10;
      q_chan1_rsci_idat_175_160 <= LOOPJ2_asn_itm_52;
      q_chan1_rsci_idat_863_848 <= LOOPJ2_asn_itm_9;
      q_chan1_rsci_idat_159_144 <= LOOPJ2_asn_itm_53;
      q_chan1_rsci_idat_879_864 <= LOOPJ2_asn_itm_8;
      q_chan1_rsci_idat_143_128 <= LOOPJ2_asn_itm_54;
      q_chan1_rsci_idat_895_880 <= LOOPJ2_asn_itm_7;
      q_chan1_rsci_idat_127_112 <= LOOPJ2_asn_itm_55;
      q_chan1_rsci_idat_911_896 <= LOOPJ2_asn_itm_6;
      q_chan1_rsci_idat_111_96 <= LOOPJ2_asn_itm_56;
      q_chan1_rsci_idat_927_912 <= LOOPJ2_asn_itm_5;
      q_chan1_rsci_idat_95_80 <= LOOPJ2_asn_itm_57;
      q_chan1_rsci_idat_943_928 <= LOOPJ2_asn_itm_4;
      q_chan1_rsci_idat_79_64 <= LOOPJ2_asn_itm_58;
      q_chan1_rsci_idat_959_944 <= LOOPJ2_asn_itm_3;
      q_chan1_rsci_idat_63_48 <= LOOPJ2_asn_itm_59;
      q_chan1_rsci_idat_975_960 <= LOOPJ2_asn_itm_2;
      q_chan1_rsci_idat_47_32 <= LOOPJ2_asn_itm_60;
      q_chan1_rsci_idat_991_976 <= LOOPJ2_asn_itm_1;
      q_chan1_rsci_idat_31_16 <= LOOPJ2_asn_itm_61;
      q_chan1_rsci_idat_1007_992 <= LOOPJ2_asn_itm;
      q_chan1_rsci_idat_15_0 <= LOOPJ2_asn_itm_62;
      q_chan1_rsci_idat_1023_1008 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_122))
        ) begin
      channel_in_data_63_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_122))
        ) begin
      channel_in_data_62_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_130))
        ) begin
      channel_in_data_1_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_122))
        ) begin
      channel_in_data_61_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_130))
        ) begin
      channel_in_data_2_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_122))
        ) begin
      channel_in_data_60_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_130))
        ) begin
      channel_in_data_3_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_122))
        ) begin
      channel_in_data_59_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_130))
        ) begin
      channel_in_data_4_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_122))
        ) begin
      channel_in_data_58_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_130))
        ) begin
      channel_in_data_5_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_122))
        ) begin
      channel_in_data_57_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_130))
        ) begin
      channel_in_data_6_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_4 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_122))
        ) begin
      channel_in_data_56_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_12 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_130))
        ) begin
      channel_in_data_7_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_153))
        ) begin
      channel_in_data_55_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_156))
        ) begin
      channel_in_data_8_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_153))
        ) begin
      channel_in_data_54_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_156))
        ) begin
      channel_in_data_9_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_153))
        ) begin
      channel_in_data_53_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_156))
        ) begin
      channel_in_data_10_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_153))
        ) begin
      channel_in_data_52_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_156))
        ) begin
      channel_in_data_11_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_153))
        ) begin
      channel_in_data_51_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_156))
        ) begin
      channel_in_data_12_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_153))
        ) begin
      channel_in_data_50_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_156))
        ) begin
      channel_in_data_13_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_153))
        ) begin
      channel_in_data_49_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_156))
        ) begin
      channel_in_data_14_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_34 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_153))
        ) begin
      channel_in_data_48_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_37 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_156))
        ) begin
      channel_in_data_15_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_172))
        ) begin
      channel_in_data_47_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_174))
        ) begin
      channel_in_data_16_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_172))
        ) begin
      channel_in_data_46_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_174))
        ) begin
      channel_in_data_17_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_172))
        ) begin
      channel_in_data_45_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_174))
        ) begin
      channel_in_data_18_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_172))
        ) begin
      channel_in_data_44_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_174))
        ) begin
      channel_in_data_19_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_172))
        ) begin
      channel_in_data_43_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_174))
        ) begin
      channel_in_data_20_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_172))
        ) begin
      channel_in_data_42_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_174))
        ) begin
      channel_in_data_21_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_172))
        ) begin
      channel_in_data_41_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_174))
        ) begin
      channel_in_data_22_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_53 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_172))
        ) begin
      channel_in_data_40_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_55 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_174))
        ) begin
      channel_in_data_23_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_190))
        ) begin
      channel_in_data_39_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_192))
        ) begin
      channel_in_data_24_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_190))
        ) begin
      channel_in_data_38_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_192))
        ) begin
      channel_in_data_25_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_190))
        ) begin
      channel_in_data_37_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_192))
        ) begin
      channel_in_data_26_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_190))
        ) begin
      channel_in_data_36_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_192))
        ) begin
      channel_in_data_27_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_22) & (~(or_dcpl_141 | or_dcpl_190))
        ) begin
      channel_in_data_35_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_20) & (~(or_dcpl_139 | or_dcpl_192))
        ) begin
      channel_in_data_28_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_18) & (~(or_dcpl_136 | or_dcpl_190))
        ) begin
      channel_in_data_34_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_15) & (~(or_dcpl_134 | or_dcpl_192))
        ) begin
      channel_in_data_29_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_9) & (~(or_dcpl_132 | or_dcpl_190))
        ) begin
      channel_in_data_33_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_6) & (~(or_dcpl_127 | or_dcpl_192))
        ) begin
      channel_in_data_30_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_71 | or_dcpl_30) & (~(or_dcpl_149 | or_dcpl_190))
        ) begin
      channel_in_data_32_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( channel_in_data_and_cse & (or_dcpl_73 | or_dcpl_1) & (~(or_dcpl_124 | or_dcpl_192))
        ) begin
      channel_in_data_31_lpi_4 <= din_chan_rsci_idat_mxwt;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_din_chan_rsci_oswt_cse <= 1'b0;
      reg_q_chan1_rsci_oswt_cse <= 1'b0;
      reg_k_chan1_rsci_oswt_cse <= 1'b0;
      reg_v_chan1_rsci_oswt_cse <= 1'b0;
      reg_pp_buf_data_rsci_oswt_1_cse <= 1'b0;
    end
    else if ( rst ) begin
      reg_din_chan_rsci_oswt_cse <= 1'b0;
      reg_q_chan1_rsci_oswt_cse <= 1'b0;
      reg_k_chan1_rsci_oswt_cse <= 1'b0;
      reg_v_chan1_rsci_oswt_cse <= 1'b0;
      reg_pp_buf_data_rsci_oswt_1_cse <= 1'b0;
    end
    else if ( run_wen ) begin
      reg_din_chan_rsci_oswt_cse <= ~(mux_57_nl | (fsm_output[7]) | (fsm_output[2])
          | or_145_cse);
      reg_q_chan1_rsci_oswt_cse <= and_dcpl_36 & and_dcpl_16 & and_dcpl_33;
      reg_k_chan1_rsci_oswt_cse <= and_dcpl_40 & and_dcpl_35 & and_dcpl_33;
      reg_v_chan1_rsci_oswt_cse <= and_dcpl_18 & and_237_cse & and_dcpl_33;
      reg_pp_buf_data_rsci_oswt_1_cse <= ~ mux_69_itm;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (and_dcpl_34 | and_dcpl_151) & ((~(or_dcpl_149 | or_dcpl_130))
        | and_dcpl_151) ) begin
      LOOPJ2_asn_itm <= MUX_v_16_2_2(din_chan_rsci_idat_mxwt, pp_buf_data_rsci_q_d_mxwt,
          and_dcpl_151);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_220)) ) begin
      LOOPJ2_asn_itm_62 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_222)) ) begin
      LOOPJ2_asn_itm_61 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_220)) ) begin
      LOOPJ2_asn_itm_60 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_222)) ) begin
      LOOPJ2_asn_itm_59 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_227)) ) begin
      LOOPJ2_asn_itm_58 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_230)) ) begin
      LOOPJ2_asn_itm_57 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_227)) ) begin
      LOOPJ2_asn_itm_56 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_230)) ) begin
      LOOPJ2_asn_itm_55 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_97 | or_dcpl_236)) ) begin
      LOOPJ2_asn_itm_54 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_97 | or_dcpl_239)) ) begin
      LOOPJ2_asn_itm_53 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_98 | or_dcpl_236)) ) begin
      LOOPJ2_asn_itm_52 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_98 | or_dcpl_239)) ) begin
      LOOPJ2_asn_itm_51 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_244)) ) begin
      LOOPJ2_asn_itm_50 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_246)) ) begin
      LOOPJ2_asn_itm_49 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_244)) ) begin
      LOOPJ2_asn_itm_48 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_246)) ) begin
      LOOPJ2_asn_itm_47 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_251)) ) begin
      LOOPJ2_asn_itm_46 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_253)) ) begin
      LOOPJ2_asn_itm_45 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_251)) ) begin
      LOOPJ2_asn_itm_44 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_253)) ) begin
      LOOPJ2_asn_itm_43 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_258)) ) begin
      LOOPJ2_asn_itm_42 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_260)) ) begin
      LOOPJ2_asn_itm_41 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_258)) ) begin
      LOOPJ2_asn_itm_40 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_260)) ) begin
      LOOPJ2_asn_itm_39 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_99 | or_dcpl_235)) ) begin
      LOOPJ2_asn_itm_38 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_99 | or_dcpl_238)) ) begin
      LOOPJ2_asn_itm_37 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_100 | or_dcpl_235)) ) begin
      LOOPJ2_asn_itm_36 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_100 | or_dcpl_238)) ) begin
      LOOPJ2_asn_itm_35 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_269)) ) begin
      LOOPJ2_asn_itm_34 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_272)) ) begin
      LOOPJ2_asn_itm_33 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_269)) ) begin
      LOOPJ2_asn_itm_32 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_272)) ) begin
      LOOPJ2_asn_itm_31 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_276)) ) begin
      LOOPJ2_asn_itm_30 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_278)) ) begin
      LOOPJ2_asn_itm_29 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_276)) ) begin
      LOOPJ2_asn_itm_28 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_278)) ) begin
      LOOPJ2_asn_itm_27 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_282)) ) begin
      LOOPJ2_asn_itm_26 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_284)) ) begin
      LOOPJ2_asn_itm_25 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_282)) ) begin
      LOOPJ2_asn_itm_24 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_284)) ) begin
      LOOPJ2_asn_itm_23 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_97 | or_dcpl_288)) ) begin
      LOOPJ2_asn_itm_22 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_97 | or_dcpl_290)) ) begin
      LOOPJ2_asn_itm_21 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_98 | or_dcpl_288)) ) begin
      LOOPJ2_asn_itm_20 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_98 | or_dcpl_290)) ) begin
      LOOPJ2_asn_itm_19 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_294)) ) begin
      LOOPJ2_asn_itm_18 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_296)) ) begin
      LOOPJ2_asn_itm_17 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_294)) ) begin
      LOOPJ2_asn_itm_16 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_296)) ) begin
      LOOPJ2_asn_itm_15 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_300)) ) begin
      LOOPJ2_asn_itm_14 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_91 | or_dcpl_302)) ) begin
      LOOPJ2_asn_itm_13 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_300)) ) begin
      LOOPJ2_asn_itm_12 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_93 | or_dcpl_302)) ) begin
      LOOPJ2_asn_itm_11 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_306)) ) begin
      LOOPJ2_asn_itm_10 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_228 | or_dcpl_308)) ) begin
      LOOPJ2_asn_itm_9 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_306)) ) begin
      LOOPJ2_asn_itm_8 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_dcpl_232 | or_dcpl_308)) ) begin
      LOOPJ2_asn_itm_7 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & nor_53_cse ) begin
      LOOPJ2_asn_itm_6 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_102 | (~ (fsm_output[0])))) ) begin
      LOOPJ2_asn_itm_5 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & nor_54_cse ) begin
      LOOPJ2_asn_itm_4 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_104 | (~ (fsm_output[0])))) ) begin
      LOOPJ2_asn_itm_3 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_106 | or_108_cse | or_dcpl_93)) ) begin
      LOOPJ2_asn_itm_2 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(mux_tmp_106 | or_dcpl_101)) ) begin
      LOOPJ2_asn_itm_1 <= pp_buf_data_rsci_q_d_mxwt;
    end
  end
  always @(posedge clk) begin
    if ( mux_162_nl & run_wen ) begin
      LOOPK2_acc_1_itm <= MUX_v_6_2_2(6'b000000, LOOPJ2_j_LOOPJ2_j_mux_nl, LOOPK2_not_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm <= 1'b0;
    end
    else if ( rst ) begin
      LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm <= 1'b0;
    end
    else if ( run_wen & (~(or_472_cse | (~ (fsm_output[2])) | ((fsm_output[6]) ^
        (fsm_output[1])) | or_dcpl_101)) ) begin
      LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm <= ~((LOOPK2_acc_1_itm != (z_out_1[5:0]))
          | (z_out_1[6]));
    end
  end
  always @(posedge clk) begin
    if ( run_wen & mux_155_nl ) begin
      LOOPK3_acc_1_itm <= z_out;
    end
  end
  always @(posedge clk) begin
    if ( LOOPJ1_j_and_ssc ) begin
      LOOPJ1_j_sva_7 <= LOOPJ1_acc_itm_7 & (~ LOOPJ1_j_sva_mx0c2);
      LOOPJ1_j_sva_6 <= (LOOPJ1_acc_itm_6_0[6]) & (~ LOOPJ1_j_sva_mx0c2);
    end
  end
  always @(posedge clk) begin
    if ( mux_165_nl & (~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[7]))) &
        (~ (fsm_output[5])) & run_wen ) begin
      LOOPJ1_j_sva_5_0 <= MUX_v_6_2_2(6'b000000, LOOPJ1_mux_65_nl, nor_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPJ1_acc_itm_7 <= 1'b0;
    end
    else if ( rst ) begin
      LOOPJ1_acc_itm_7 <= 1'b0;
    end
    else if ( run_wen & ((~ mux_125_nl) | and_dcpl_153) ) begin
      LOOPJ1_acc_itm_7 <= LOOPJ1_acc_sdt[7];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOPJ1_acc_itm_6_0 <= 7'b0000000;
    end
    else if ( rst ) begin
      LOOPJ1_acc_itm_6_0 <= 7'b0000000;
    end
    else if ( mux_169_nl & nor_145_cse & run_wen ) begin
      LOOPJ1_acc_itm_6_0 <= MUX_v_7_2_2(LOOPK1_k_and_nl, (LOOPJ1_acc_sdt[6:0]), and_dcpl_153);
    end
  end
  assign LOOPI1_i_not_1_nl = ~ LOOPI1_i_sva_mx0c0;
  assign mux_54_nl = MUX_s_1_2_2(mux_tmp_53, or_tmp_46, fsm_output[3]);
  assign or_259_nl = (fsm_output[3]) | mux_tmp_53;
  assign mux_55_nl = MUX_s_1_2_2(mux_54_nl, or_259_nl, LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp);
  assign or_258_nl = (fsm_output[1]) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_51_nl = MUX_s_1_2_2(or_258_nl, or_tmp_46, fsm_output[3]);
  assign or_255_nl = (fsm_output[3]) | (fsm_output[1]) | (fsm_output[6]) | (fsm_output[8]);
  assign mux_52_nl = MUX_s_1_2_2(mux_51_nl, or_255_nl, LOOPI1_LOOPI1_if_LOOPI1_if_nor_tmp);
  assign mux_56_nl = MUX_s_1_2_2(mux_55_nl, mux_52_nl, LOOPJ1_LOOPJ1_if_LOOPJ1_if_nor_tmp);
  assign or_254_nl = LOOPK1_LOOPK1_if_1_LOOPK1_if_1_nor_tmp | (fsm_output[3]) | (fsm_output[1])
      | (fsm_output[6]) | (fsm_output[8]);
  assign mux_57_nl = MUX_s_1_2_2(mux_56_nl, or_254_nl, fsm_output[0]);
  assign and_223_nl = and_dcpl_18 & and_dcpl_9 & and_dcpl_15;
  assign LOOPJ2_j_LOOPJ2_j_mux_nl = MUX_v_6_2_2(z_out, LOOPK3_acc_1_itm, and_223_nl);
  assign or_452_nl = ((fsm_output[6]) & LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm) | (fsm_output[8:7]!=2'b01);
  assign mux_144_nl = MUX_s_1_2_2(mux_tmp_143, or_452_nl, fsm_output[1]);
  assign or_451_nl = (fsm_output[1]) | (fsm_output[6]);
  assign mux_142_nl = MUX_s_1_2_2(mux_tmp_140, or_472_cse, or_451_nl);
  assign mux_145_nl = MUX_s_1_2_2(mux_144_nl, mux_142_nl, fsm_output[0]);
  assign mux_146_nl = MUX_s_1_2_2(mux_tmp_143, mux_145_nl, fsm_output[2]);
  assign or_450_nl = (fsm_output[2]) | (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]);
  assign mux_141_nl = MUX_s_1_2_2(mux_tmp_140, or_472_cse, or_450_nl);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, mux_141_nl, fsm_output[3]);
  assign mux_148_nl = MUX_s_1_2_2(mux_147_nl, or_472_cse, or_145_cse);
  assign LOOPK2_not_nl = ~ mux_148_nl;
  assign mux_160_nl = MUX_s_1_2_2(or_478_cse, or_146_cse_1, fsm_output[7]);
  assign mux_nl = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), fsm_output[1]);
  assign nor_135_nl = ~((fsm_output[1]) | (fsm_output[6]));
  assign or_473_nl = (~ LOOPK2_LOOPK2_if_LOOPK2_if_nor_itm) | (fsm_output[0]);
  assign mux_158_nl = MUX_s_1_2_2(mux_nl, nor_135_nl, or_473_nl);
  assign or_475_nl = (fsm_output[8]) | mux_158_nl;
  assign mux_159_nl = MUX_s_1_2_2(or_476_cse, or_475_nl, fsm_output[7]);
  assign mux_161_nl = MUX_s_1_2_2(mux_160_nl, mux_159_nl, fsm_output[2]);
  assign mux_162_nl = MUX_s_1_2_2(mux_161_nl, or_472_cse, or_158_cse_1);
  assign mux_155_nl = MUX_s_1_2_2(or_dcpl_104, or_dcpl_109, or_158_cse_1);
  assign LOOPJ1_mux_65_nl = MUX_v_6_2_2(z_out, (LOOPJ1_acc_itm_6_0[5:0]), mux_36_itm);
  assign mux_170_nl = MUX_s_1_2_2(mux_tmp_34, mux_tmp_31, fsm_output[0]);
  assign mux_171_nl = MUX_s_1_2_2(mux_170_nl, or_tmp_23, fsm_output[5]);
  assign nor_nl = ~((mux_171_nl & (~ mux_36_itm)) | LOOPJ1_j_sva_mx0c2);
  assign nor_136_nl = ~((fsm_output[0]) | (fsm_output[3]) | (fsm_output[1]));
  assign nor_137_nl = ~((fsm_output[0]) | (fsm_output[3]) | (~ (fsm_output[1])));
  assign mux_164_nl = MUX_s_1_2_2(nor_136_nl, nor_137_nl, fsm_output[6]);
  assign nand_27_nl = ~((fsm_output[3]) & (fsm_output[1]));
  assign or_479_nl = (~ (fsm_output[3])) | (fsm_output[1]);
  assign mux_163_nl = MUX_s_1_2_2(nand_27_nl, or_479_nl, fsm_output[0]);
  assign nor_138_nl = ~((fsm_output[6]) | mux_163_nl);
  assign mux_165_nl = MUX_s_1_2_2(mux_164_nl, nor_138_nl, fsm_output[8]);
  assign nor_55_nl = ~((~ (fsm_output[1])) | (fsm_output[8]));
  assign or_346_nl = (fsm_output[0]) | (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_121_nl = MUX_s_1_2_2(nor_55_nl, or_346_nl, fsm_output[6]);
  assign mux_122_nl = MUX_s_1_2_2(mux_121_nl, or_146_cse_1, fsm_output[7]);
  assign or_344_nl = (fsm_output[6]) | (fsm_output[0]) | (~((fsm_output[1]) & (fsm_output[8])));
  assign mux_129_nl = MUX_s_1_2_2(or_344_nl, (fsm_output[8]), fsm_output[7]);
  assign mux_123_nl = MUX_s_1_2_2(mux_122_nl, mux_129_nl, fsm_output[3]);
  assign or_340_nl = nor_49_cse | (fsm_output[8]);
  assign or_326_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[8]);
  assign mux_126_nl = MUX_s_1_2_2(or_340_nl, or_326_nl, fsm_output[6]);
  assign mux_127_nl = MUX_s_1_2_2(or_476_cse, mux_126_nl, fsm_output[7]);
  assign mux_128_nl = MUX_s_1_2_2(mux_127_nl, or_472_cse, fsm_output[3]);
  assign mux_124_nl = MUX_s_1_2_2(mux_123_nl, mux_128_nl, fsm_output[2]);
  assign mux_125_nl = MUX_s_1_2_2(mux_124_nl, or_472_cse, or_145_cse);
  assign LOOPK1_k_mux1h_nl = MUX1HOT_v_7_3_2(LOOPK1_acc_1_tmp, LOOPK2_acc_tmp_sva_mx0w2,
      LOOPK3_acc_psp_sva_mx0w4, {and_dcpl_34 , and_dcpl_38 , and_dcpl_42});
  assign nor_59_nl = ~((fsm_output[6:0]!=7'b0000001));
  assign or_466_nl = (((fsm_output[1:0]!=2'b00)) & (fsm_output[2])) | (fsm_output[5:3]!=3'b000);
  assign or_467_nl = ((fsm_output[1:0]==2'b11)) | (fsm_output[5:2]!=4'b0001);
  assign mux_43_nl = MUX_s_1_2_2(or_466_nl, or_467_nl, fsm_output[6]);
  assign mux_44_nl = MUX_s_1_2_2(nor_59_nl, mux_43_nl, fsm_output[7]);
  assign nor_60_nl = ~((fsm_output[7:6]!=2'b00) | and_237_cse | (fsm_output[5:3]!=3'b000));
  assign mux_45_nl = MUX_s_1_2_2(mux_44_nl, nor_60_nl, fsm_output[8]);
  assign LOOPK1_k_and_nl = MUX_v_7_2_2(7'b0000000, LOOPK1_k_mux1h_nl, mux_45_nl);
  assign nor_141_nl = ~((fsm_output[3]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[8]));
  assign nor_142_nl = ~((~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[2]))
      | (fsm_output[6]) | (fsm_output[8]));
  assign mux_168_nl = MUX_s_1_2_2(nor_141_nl, nor_142_nl, fsm_output[7]);
  assign or_487_nl = (fsm_output[2]) | (fsm_output[8]);
  assign or_486_nl = (fsm_output[2]) | (fsm_output[6]) | (~ (fsm_output[8]));
  assign mux_166_nl = MUX_s_1_2_2(or_487_nl, or_486_nl, fsm_output[3]);
  assign nor_143_nl = ~((fsm_output[0]) | mux_166_nl);
  assign nor_144_nl = ~((~ (fsm_output[0])) | (fsm_output[3]) | (~ (fsm_output[2]))
      | (~ (fsm_output[6])) | (fsm_output[8]));
  assign mux_167_nl = MUX_s_1_2_2(nor_143_nl, nor_144_nl, fsm_output[7]);
  assign mux_169_nl = MUX_s_1_2_2(mux_168_nl, mux_167_nl, fsm_output[1]);
  assign LOOPI1_mux_1_nl = MUX_v_2_2_2((LOOPK2_acc_1_itm[5:4]), (LOOPJ1_j_sva_5_0[5:4]),
      and_263_itm);
  assign not_457_nl = ~ and_252_itm;
  assign LOOPI1_LOOPI1_and_1_nl = MUX_v_2_2_2(2'b00, LOOPI1_mux_1_nl, not_457_nl);
  assign and_301_nl = nor_145_cse & (~ (fsm_output[3])) & (~((fsm_output[1]) ^ (fsm_output[6])))
      & (fsm_output[2]) & (fsm_output[0]) & (fsm_output[7]) & (~ (fsm_output[8]));
  assign LOOPI1_mux1h_2_nl = MUX1HOT_v_4_3_2(LOOPI1_i_sva, (LOOPK2_acc_1_itm[3:0]),
      (LOOPJ1_j_sva_5_0[3:0]), {and_252_itm , and_301_nl , and_263_itm});
  assign nl_z_out = ({LOOPI1_LOOPI1_and_1_nl , LOOPI1_mux1h_2_nl}) + 6'b000001;
  assign z_out = nl_z_out[5:0];
  assign operator_7_false_operator_7_false_and_2_nl = (dim[6]) & (~(and_277_itm |
      and_280_itm | and_286_itm));
  assign operator_7_false_mux_1_nl = MUX_s_1_2_2((dim[5]), (length[5]), and_280_itm);
  assign operator_7_false_operator_7_false_and_3_nl = operator_7_false_mux_1_nl &
      (~(and_277_itm | and_286_itm));
  assign operator_7_false_mux1h_4_nl = MUX1HOT_s_1_3_2((dim[4]), (length[5]), (length[4]),
      {and_271_itm , and_277_itm , and_280_itm});
  assign operator_7_false_and_1_nl = operator_7_false_mux1h_4_nl & (~ and_286_itm);
  assign operator_7_false_mux1h_5_nl = MUX1HOT_v_4_4_2((dim[3:0]), (length[4:1]),
      (length[3:0]), head, {and_271_itm , and_277_itm , and_280_itm , and_286_itm});
  assign nl_z_out_1 = conv_u2u_7_8({operator_7_false_operator_7_false_and_2_nl ,
      operator_7_false_operator_7_false_and_3_nl , operator_7_false_and_1_nl , operator_7_false_mux1h_5_nl})
      + 8'b11111111;
  assign z_out_1 = nl_z_out_1[7:0];

  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [15:0] MUX1HOT_v_16_64_2;
    input [15:0] input_63;
    input [15:0] input_62;
    input [15:0] input_61;
    input [15:0] input_60;
    input [15:0] input_59;
    input [15:0] input_58;
    input [15:0] input_57;
    input [15:0] input_56;
    input [15:0] input_55;
    input [15:0] input_54;
    input [15:0] input_53;
    input [15:0] input_52;
    input [15:0] input_51;
    input [15:0] input_50;
    input [15:0] input_49;
    input [15:0] input_48;
    input [15:0] input_47;
    input [15:0] input_46;
    input [15:0] input_45;
    input [15:0] input_44;
    input [15:0] input_43;
    input [15:0] input_42;
    input [15:0] input_41;
    input [15:0] input_40;
    input [15:0] input_39;
    input [15:0] input_38;
    input [15:0] input_37;
    input [15:0] input_36;
    input [15:0] input_35;
    input [15:0] input_34;
    input [15:0] input_33;
    input [15:0] input_32;
    input [15:0] input_31;
    input [15:0] input_30;
    input [15:0] input_29;
    input [15:0] input_28;
    input [15:0] input_27;
    input [15:0] input_26;
    input [15:0] input_25;
    input [15:0] input_24;
    input [15:0] input_23;
    input [15:0] input_22;
    input [15:0] input_21;
    input [15:0] input_20;
    input [15:0] input_19;
    input [15:0] input_18;
    input [15:0] input_17;
    input [15:0] input_16;
    input [15:0] input_15;
    input [15:0] input_14;
    input [15:0] input_13;
    input [15:0] input_12;
    input [15:0] input_11;
    input [15:0] input_10;
    input [15:0] input_9;
    input [15:0] input_8;
    input [15:0] input_7;
    input [15:0] input_6;
    input [15:0] input_5;
    input [15:0] input_4;
    input [15:0] input_3;
    input [15:0] input_2;
    input [15:0] input_1;
    input [15:0] input_0;
    input [63:0] sel;
    reg [15:0] result;
  begin
    result = input_0 & {16{sel[0]}};
    result = result | (input_1 & {16{sel[1]}});
    result = result | (input_2 & {16{sel[2]}});
    result = result | (input_3 & {16{sel[3]}});
    result = result | (input_4 & {16{sel[4]}});
    result = result | (input_5 & {16{sel[5]}});
    result = result | (input_6 & {16{sel[6]}});
    result = result | (input_7 & {16{sel[7]}});
    result = result | (input_8 & {16{sel[8]}});
    result = result | (input_9 & {16{sel[9]}});
    result = result | (input_10 & {16{sel[10]}});
    result = result | (input_11 & {16{sel[11]}});
    result = result | (input_12 & {16{sel[12]}});
    result = result | (input_13 & {16{sel[13]}});
    result = result | (input_14 & {16{sel[14]}});
    result = result | (input_15 & {16{sel[15]}});
    result = result | (input_16 & {16{sel[16]}});
    result = result | (input_17 & {16{sel[17]}});
    result = result | (input_18 & {16{sel[18]}});
    result = result | (input_19 & {16{sel[19]}});
    result = result | (input_20 & {16{sel[20]}});
    result = result | (input_21 & {16{sel[21]}});
    result = result | (input_22 & {16{sel[22]}});
    result = result | (input_23 & {16{sel[23]}});
    result = result | (input_24 & {16{sel[24]}});
    result = result | (input_25 & {16{sel[25]}});
    result = result | (input_26 & {16{sel[26]}});
    result = result | (input_27 & {16{sel[27]}});
    result = result | (input_28 & {16{sel[28]}});
    result = result | (input_29 & {16{sel[29]}});
    result = result | (input_30 & {16{sel[30]}});
    result = result | (input_31 & {16{sel[31]}});
    result = result | (input_32 & {16{sel[32]}});
    result = result | (input_33 & {16{sel[33]}});
    result = result | (input_34 & {16{sel[34]}});
    result = result | (input_35 & {16{sel[35]}});
    result = result | (input_36 & {16{sel[36]}});
    result = result | (input_37 & {16{sel[37]}});
    result = result | (input_38 & {16{sel[38]}});
    result = result | (input_39 & {16{sel[39]}});
    result = result | (input_40 & {16{sel[40]}});
    result = result | (input_41 & {16{sel[41]}});
    result = result | (input_42 & {16{sel[42]}});
    result = result | (input_43 & {16{sel[43]}});
    result = result | (input_44 & {16{sel[44]}});
    result = result | (input_45 & {16{sel[45]}});
    result = result | (input_46 & {16{sel[46]}});
    result = result | (input_47 & {16{sel[47]}});
    result = result | (input_48 & {16{sel[48]}});
    result = result | (input_49 & {16{sel[49]}});
    result = result | (input_50 & {16{sel[50]}});
    result = result | (input_51 & {16{sel[51]}});
    result = result | (input_52 & {16{sel[52]}});
    result = result | (input_53 & {16{sel[53]}});
    result = result | (input_54 & {16{sel[54]}});
    result = result | (input_55 & {16{sel[55]}});
    result = result | (input_56 & {16{sel[56]}});
    result = result | (input_57 & {16{sel[57]}});
    result = result | (input_58 & {16{sel[58]}});
    result = result | (input_59 & {16{sel[59]}});
    result = result | (input_60 & {16{sel[60]}});
    result = result | (input_61 & {16{sel[61]}});
    result = result | (input_62 & {16{sel[62]}});
    result = result | (input_63 & {16{sel[63]}});
    MUX1HOT_v_16_64_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_62_2;
    input [5:0] input_61;
    input [5:0] input_60;
    input [5:0] input_59;
    input [5:0] input_58;
    input [5:0] input_57;
    input [5:0] input_56;
    input [5:0] input_55;
    input [5:0] input_54;
    input [5:0] input_53;
    input [5:0] input_52;
    input [5:0] input_51;
    input [5:0] input_50;
    input [5:0] input_49;
    input [5:0] input_48;
    input [5:0] input_47;
    input [5:0] input_46;
    input [5:0] input_45;
    input [5:0] input_44;
    input [5:0] input_43;
    input [5:0] input_42;
    input [5:0] input_41;
    input [5:0] input_40;
    input [5:0] input_39;
    input [5:0] input_38;
    input [5:0] input_37;
    input [5:0] input_36;
    input [5:0] input_35;
    input [5:0] input_34;
    input [5:0] input_33;
    input [5:0] input_32;
    input [5:0] input_31;
    input [5:0] input_30;
    input [5:0] input_29;
    input [5:0] input_28;
    input [5:0] input_27;
    input [5:0] input_26;
    input [5:0] input_25;
    input [5:0] input_24;
    input [5:0] input_23;
    input [5:0] input_22;
    input [5:0] input_21;
    input [5:0] input_20;
    input [5:0] input_19;
    input [5:0] input_18;
    input [5:0] input_17;
    input [5:0] input_16;
    input [5:0] input_15;
    input [5:0] input_14;
    input [5:0] input_13;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [61:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    result = result | (input_9 & {6{sel[9]}});
    result = result | (input_10 & {6{sel[10]}});
    result = result | (input_11 & {6{sel[11]}});
    result = result | (input_12 & {6{sel[12]}});
    result = result | (input_13 & {6{sel[13]}});
    result = result | (input_14 & {6{sel[14]}});
    result = result | (input_15 & {6{sel[15]}});
    result = result | (input_16 & {6{sel[16]}});
    result = result | (input_17 & {6{sel[17]}});
    result = result | (input_18 & {6{sel[18]}});
    result = result | (input_19 & {6{sel[19]}});
    result = result | (input_20 & {6{sel[20]}});
    result = result | (input_21 & {6{sel[21]}});
    result = result | (input_22 & {6{sel[22]}});
    result = result | (input_23 & {6{sel[23]}});
    result = result | (input_24 & {6{sel[24]}});
    result = result | (input_25 & {6{sel[25]}});
    result = result | (input_26 & {6{sel[26]}});
    result = result | (input_27 & {6{sel[27]}});
    result = result | (input_28 & {6{sel[28]}});
    result = result | (input_29 & {6{sel[29]}});
    result = result | (input_30 & {6{sel[30]}});
    result = result | (input_31 & {6{sel[31]}});
    result = result | (input_32 & {6{sel[32]}});
    result = result | (input_33 & {6{sel[33]}});
    result = result | (input_34 & {6{sel[34]}});
    result = result | (input_35 & {6{sel[35]}});
    result = result | (input_36 & {6{sel[36]}});
    result = result | (input_37 & {6{sel[37]}});
    result = result | (input_38 & {6{sel[38]}});
    result = result | (input_39 & {6{sel[39]}});
    result = result | (input_40 & {6{sel[40]}});
    result = result | (input_41 & {6{sel[41]}});
    result = result | (input_42 & {6{sel[42]}});
    result = result | (input_43 & {6{sel[43]}});
    result = result | (input_44 & {6{sel[44]}});
    result = result | (input_45 & {6{sel[45]}});
    result = result | (input_46 & {6{sel[46]}});
    result = result | (input_47 & {6{sel[47]}});
    result = result | (input_48 & {6{sel[48]}});
    result = result | (input_49 & {6{sel[49]}});
    result = result | (input_50 & {6{sel[50]}});
    result = result | (input_51 & {6{sel[51]}});
    result = result | (input_52 & {6{sel[52]}});
    result = result | (input_53 & {6{sel[53]}});
    result = result | (input_54 & {6{sel[54]}});
    result = result | (input_55 & {6{sel[55]}});
    result = result | (input_56 & {6{sel[56]}});
    result = result | (input_57 & {6{sel[57]}});
    result = result | (input_58 & {6{sel[58]}});
    result = result | (input_59 & {6{sel[59]}});
    result = result | (input_60 & {6{sel[60]}});
    result = result | (input_61 & {6{sel[61]}});
    MUX1HOT_v_6_62_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input  sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [8:0] conv_s2s_7_9 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_9 = {{2{vector[6]}}, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_7_9 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_9 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2u_5_7 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_7 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Buffer
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Buffer (
  clk, rst, arst_n, head, length, dim, din_chan_rsc_dat, din_chan_rsc_vld, din_chan_rsc_rdy,
      q_chan1_rsc_dat, q_chan1_rsc_vld, q_chan1_rsc_rdy, k_chan1_rsc_dat, k_chan1_rsc_vld,
      k_chan1_rsc_rdy, v_chan1_rsc_dat, v_chan1_rsc_vld, v_chan1_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [15:0] din_chan_rsc_dat;
  input din_chan_rsc_vld;
  output din_chan_rsc_rdy;
  output [1023:0] q_chan1_rsc_dat;
  output q_chan1_rsc_vld;
  input q_chan1_rsc_rdy;
  output [1023:0] k_chan1_rsc_dat;
  output k_chan1_rsc_vld;
  input k_chan1_rsc_rdy;
  output [1023:0] v_chan1_rsc_dat;
  output v_chan1_rsc_vld;
  input v_chan1_rsc_rdy;


  // Interconnect Declarations
  wire [13:0] pp_buf_data_rsci_radr_d;
  wire [13:0] pp_buf_data_rsci_wadr_d;
  wire [15:0] pp_buf_data_rsci_d_d;
  wire [15:0] pp_buf_data_rsci_q_d;
  wire pp_buf_data_rsc_we;
  wire [15:0] pp_buf_data_rsc_d;
  wire [13:0] pp_buf_data_rsc_wadr;
  wire [15:0] pp_buf_data_rsc_q;
  wire pp_buf_data_rsc_re;
  wire [13:0] pp_buf_data_rsc_radr;
  wire pp_buf_data_rsci_we_d_iff;
  wire pp_buf_data_rsci_re_d_iff;


  // Interconnect Declarations for Component Instantiations 
  ccs_ram_sync_1R1W #(.data_width(32'sd16),
  .addr_width(32'sd14),
  .depth(32'sd10752)) pp_buf_data_rsc_comp (
      .radr(pp_buf_data_rsc_radr),
      .wadr(pp_buf_data_rsc_wadr),
      .d(pp_buf_data_rsc_d),
      .we(pp_buf_data_rsc_we),
      .re(pp_buf_data_rsc_re),
      .clk(clk),
      .q(pp_buf_data_rsc_q)
    );
  ATTENTION_IP_Attention_Buffer_ccs_sample_mem_ccs_ram_sync_1R1W_rwport_8_16_14_10752_10752_16_5_gen
      pp_buf_data_rsci (
      .we(pp_buf_data_rsc_we),
      .d(pp_buf_data_rsc_d),
      .wadr(pp_buf_data_rsc_wadr),
      .q(pp_buf_data_rsc_q),
      .re(pp_buf_data_rsc_re),
      .radr(pp_buf_data_rsc_radr),
      .radr_d(pp_buf_data_rsci_radr_d),
      .wadr_d(pp_buf_data_rsci_wadr_d),
      .d_d(pp_buf_data_rsci_d_d),
      .we_d(pp_buf_data_rsci_we_d_iff),
      .re_d(pp_buf_data_rsci_re_d_iff),
      .q_d(pp_buf_data_rsci_q_d),
      .port_0_r_ram_ir_internal_RMASK_B_d(pp_buf_data_rsci_re_d_iff),
      .port_1_w_ram_ir_internal_WMASK_B_d(pp_buf_data_rsci_we_d_iff)
    );
  ATTENTION_IP_Attention_Buffer_run ATTENTION_IP_Attention_Buffer_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .din_chan_rsc_dat(din_chan_rsc_dat),
      .din_chan_rsc_vld(din_chan_rsc_vld),
      .din_chan_rsc_rdy(din_chan_rsc_rdy),
      .q_chan1_rsc_dat(q_chan1_rsc_dat),
      .q_chan1_rsc_vld(q_chan1_rsc_vld),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy),
      .k_chan1_rsc_dat(k_chan1_rsc_dat),
      .k_chan1_rsc_vld(k_chan1_rsc_vld),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy),
      .v_chan1_rsc_dat(v_chan1_rsc_dat),
      .v_chan1_rsc_vld(v_chan1_rsc_vld),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy),
      .pp_buf_data_rsci_radr_d(pp_buf_data_rsci_radr_d),
      .pp_buf_data_rsci_wadr_d(pp_buf_data_rsci_wadr_d),
      .pp_buf_data_rsci_d_d(pp_buf_data_rsci_d_d),
      .pp_buf_data_rsci_q_d(pp_buf_data_rsci_q_d),
      .pp_buf_data_rsci_we_d_pff(pp_buf_data_rsci_we_d_iff),
      .pp_buf_data_rsci_re_d_pff(pp_buf_data_rsci_re_d_iff)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   b08092@cad29.ee.ntu.edu.tw
//  Generated date: Wed Jun 12 20:45:07 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    ATTENTION_IP_Attention_Top
// ------------------------------------------------------------------


module ATTENTION_IP_Attention_Top (
  clk, rst, arst_n, head, length, dim, din_chan_rsc_dat, din_chan_rsc_vld, din_chan_rsc_rdy,
      dout_chan_rsc_dat, dout_chan_rsc_vld, dout_chan_rsc_rdy
);
  input clk;
  input rst;
  input arst_n;
  input [3:0] head;
  input [5:0] length;
  input [6:0] dim;
  input [15:0] din_chan_rsc_dat;
  input din_chan_rsc_vld;
  output din_chan_rsc_rdy;
  output [15:0] dout_chan_rsc_dat;
  output dout_chan_rsc_vld;
  input dout_chan_rsc_rdy;


  // Interconnect Declarations
  wire [1023:0] q_chan1_rsc_dat_n_Buffer_inst;
  wire [1023:0] k_chan1_rsc_dat_n_Buffer_inst;
  wire [1023:0] v_chan1_rsc_dat_n_Buffer_inst;
  wire [1023:0] q_chan2_rsc_dat_n_Filter_inst;
  wire [1023:0] k_chan2_rsc_dat_n_Filter_inst;
  wire [1023:0] v_chan2_rsc_dat_n_Filter_inst;
  wire [15:0] dout_chan_rsc_dat_n_Calculator_inst;
  wire din_chan_rsc_rdy_n_Buffer_inst_bud;
  wire q_chan1_rsc_vld_n_Buffer_inst_bud;
  wire q_chan1_rsc_rdy_n_Filter_inst_bud;
  wire k_chan1_rsc_vld_n_Buffer_inst_bud;
  wire k_chan1_rsc_rdy_n_Filter_inst_bud;
  wire v_chan1_rsc_vld_n_Buffer_inst_bud;
  wire v_chan1_rsc_rdy_n_Filter_inst_bud;
  wire q_chan2_rsc_vld_n_Filter_inst_bud;
  wire q_chan2_rsc_rdy_n_Calculator_inst_bud;
  wire k_chan2_rsc_vld_n_Filter_inst_bud;
  wire k_chan2_rsc_rdy_n_Calculator_inst_bud;
  wire v_chan2_rsc_vld_n_Filter_inst_bud;
  wire v_chan2_rsc_rdy_n_Calculator_inst_bud;
  wire dout_chan_rsc_vld_n_Calculator_inst_bud;


  // Interconnect Declarations for Component Instantiations 
  ATTENTION_IP_Attention_Buffer Buffer_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .din_chan_rsc_dat(din_chan_rsc_dat),
      .din_chan_rsc_vld(din_chan_rsc_vld),
      .din_chan_rsc_rdy(din_chan_rsc_rdy_n_Buffer_inst_bud),
      .q_chan1_rsc_dat(q_chan1_rsc_dat_n_Buffer_inst),
      .q_chan1_rsc_vld(q_chan1_rsc_vld_n_Buffer_inst_bud),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy_n_Filter_inst_bud),
      .k_chan1_rsc_dat(k_chan1_rsc_dat_n_Buffer_inst),
      .k_chan1_rsc_vld(k_chan1_rsc_vld_n_Buffer_inst_bud),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy_n_Filter_inst_bud),
      .v_chan1_rsc_dat(v_chan1_rsc_dat_n_Buffer_inst),
      .v_chan1_rsc_vld(v_chan1_rsc_vld_n_Buffer_inst_bud),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy_n_Filter_inst_bud)
    );
  ATTENTION_IP_Attention_Filter Filter_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .q_chan1_rsc_dat(q_chan1_rsc_dat_n_Buffer_inst),
      .q_chan1_rsc_vld(q_chan1_rsc_vld_n_Buffer_inst_bud),
      .q_chan1_rsc_rdy(q_chan1_rsc_rdy_n_Filter_inst_bud),
      .k_chan1_rsc_dat(k_chan1_rsc_dat_n_Buffer_inst),
      .k_chan1_rsc_vld(k_chan1_rsc_vld_n_Buffer_inst_bud),
      .k_chan1_rsc_rdy(k_chan1_rsc_rdy_n_Filter_inst_bud),
      .v_chan1_rsc_dat(v_chan1_rsc_dat_n_Buffer_inst),
      .v_chan1_rsc_vld(v_chan1_rsc_vld_n_Buffer_inst_bud),
      .v_chan1_rsc_rdy(v_chan1_rsc_rdy_n_Filter_inst_bud),
      .q_chan2_rsc_dat(q_chan2_rsc_dat_n_Filter_inst),
      .q_chan2_rsc_vld(q_chan2_rsc_vld_n_Filter_inst_bud),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy_n_Calculator_inst_bud),
      .k_chan2_rsc_dat(k_chan2_rsc_dat_n_Filter_inst),
      .k_chan2_rsc_vld(k_chan2_rsc_vld_n_Filter_inst_bud),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy_n_Calculator_inst_bud),
      .v_chan2_rsc_dat(v_chan2_rsc_dat_n_Filter_inst),
      .v_chan2_rsc_vld(v_chan2_rsc_vld_n_Filter_inst_bud),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy_n_Calculator_inst_bud)
    );
  ATTENTION_IP_Attention_Calculator Calculator_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .head(head),
      .length(length),
      .dim(dim),
      .q_chan2_rsc_dat(q_chan2_rsc_dat_n_Filter_inst),
      .q_chan2_rsc_vld(q_chan2_rsc_vld_n_Filter_inst_bud),
      .q_chan2_rsc_rdy(q_chan2_rsc_rdy_n_Calculator_inst_bud),
      .k_chan2_rsc_dat(k_chan2_rsc_dat_n_Filter_inst),
      .k_chan2_rsc_vld(k_chan2_rsc_vld_n_Filter_inst_bud),
      .k_chan2_rsc_rdy(k_chan2_rsc_rdy_n_Calculator_inst_bud),
      .v_chan2_rsc_dat(v_chan2_rsc_dat_n_Filter_inst),
      .v_chan2_rsc_vld(v_chan2_rsc_vld_n_Filter_inst_bud),
      .v_chan2_rsc_rdy(v_chan2_rsc_rdy_n_Calculator_inst_bud),
      .dout_chan_rsc_dat(dout_chan_rsc_dat_n_Calculator_inst),
      .dout_chan_rsc_vld(dout_chan_rsc_vld_n_Calculator_inst_bud),
      .dout_chan_rsc_rdy(dout_chan_rsc_rdy)
    );
  assign din_chan_rsc_rdy = din_chan_rsc_rdy_n_Buffer_inst_bud;
  assign dout_chan_rsc_vld = dout_chan_rsc_vld_n_Calculator_inst_bud;
  assign dout_chan_rsc_dat = dout_chan_rsc_dat_n_Calculator_inst;
endmodule




