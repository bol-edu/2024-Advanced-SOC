
//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld, VDD, VSS);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;
  input VDD;
  input VSS;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /usr/cadtool/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld, VDD, VSS);

  parameter integer rscid = 1;
  parameter integer width = 8;
  input VDD;
  input VSS;
  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> ./rtl_AES128_ENmgc_rom_18_256_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m112061603@ws34
//  Generated date: Sun Jun  9 02:20:57 2024
// ----------------------------------------------------------------------

// 
module AES128_ENmgc_rom_18_256_8_1 (addr, data_out, VDD, VSS
);
  input VDD;
  input VSS;
  input [7:0]addr ;
  output [7:0]data_out ;


  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 256;
  parameter n_numports = 1;
  parameter n_addr_w   = 8;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [255:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b01100011;
    mem[1] <= 8'b01111100;
    mem[2] <= 8'b01110111;
    mem[3] <= 8'b01111011;
    mem[4] <= 8'b11110010;
    mem[5] <= 8'b01101011;
    mem[6] <= 8'b01101111;
    mem[7] <= 8'b11000101;
    mem[8] <= 8'b00110000;
    mem[9] <= 8'b00000001;
    mem[10] <= 8'b01100111;
    mem[11] <= 8'b00101011;
    mem[12] <= 8'b11111110;
    mem[13] <= 8'b11010111;
    mem[14] <= 8'b10101011;
    mem[15] <= 8'b01110110;
    mem[16] <= 8'b11001010;
    mem[17] <= 8'b10000010;
    mem[18] <= 8'b11001001;
    mem[19] <= 8'b01111101;
    mem[20] <= 8'b11111010;
    mem[21] <= 8'b01011001;
    mem[22] <= 8'b01000111;
    mem[23] <= 8'b11110000;
    mem[24] <= 8'b10101101;
    mem[25] <= 8'b11010100;
    mem[26] <= 8'b10100010;
    mem[27] <= 8'b10101111;
    mem[28] <= 8'b10011100;
    mem[29] <= 8'b10100100;
    mem[30] <= 8'b01110010;
    mem[31] <= 8'b11000000;
    mem[32] <= 8'b10110111;
    mem[33] <= 8'b11111101;
    mem[34] <= 8'b10010011;
    mem[35] <= 8'b00100110;
    mem[36] <= 8'b00110110;
    mem[37] <= 8'b00111111;
    mem[38] <= 8'b11110111;
    mem[39] <= 8'b11001100;
    mem[40] <= 8'b00110100;
    mem[41] <= 8'b10100101;
    mem[42] <= 8'b11100101;
    mem[43] <= 8'b11110001;
    mem[44] <= 8'b01110001;
    mem[45] <= 8'b11011000;
    mem[46] <= 8'b00110001;
    mem[47] <= 8'b00010101;
    mem[48] <= 8'b00000100;
    mem[49] <= 8'b11000111;
    mem[50] <= 8'b00100011;
    mem[51] <= 8'b11000011;
    mem[52] <= 8'b00011000;
    mem[53] <= 8'b10010110;
    mem[54] <= 8'b00000101;
    mem[55] <= 8'b10011010;
    mem[56] <= 8'b00000111;
    mem[57] <= 8'b00010010;
    mem[58] <= 8'b10000000;
    mem[59] <= 8'b11100010;
    mem[60] <= 8'b11101011;
    mem[61] <= 8'b00100111;
    mem[62] <= 8'b10110010;
    mem[63] <= 8'b01110101;
    mem[64] <= 8'b00001001;
    mem[65] <= 8'b10000011;
    mem[66] <= 8'b00101100;
    mem[67] <= 8'b00011010;
    mem[68] <= 8'b00011011;
    mem[69] <= 8'b01101110;
    mem[70] <= 8'b01011010;
    mem[71] <= 8'b10100000;
    mem[72] <= 8'b01010010;
    mem[73] <= 8'b00111011;
    mem[74] <= 8'b11010110;
    mem[75] <= 8'b10110011;
    mem[76] <= 8'b00101001;
    mem[77] <= 8'b11100011;
    mem[78] <= 8'b00101111;
    mem[79] <= 8'b10000100;
    mem[80] <= 8'b01010011;
    mem[81] <= 8'b11010001;
    mem[82] <= 8'b00000000;
    mem[83] <= 8'b11101101;
    mem[84] <= 8'b00100000;
    mem[85] <= 8'b11111100;
    mem[86] <= 8'b10110001;
    mem[87] <= 8'b01011011;
    mem[88] <= 8'b01101010;
    mem[89] <= 8'b11001011;
    mem[90] <= 8'b10111110;
    mem[91] <= 8'b00111001;
    mem[92] <= 8'b01001010;
    mem[93] <= 8'b01001100;
    mem[94] <= 8'b01011000;
    mem[95] <= 8'b11001111;
    mem[96] <= 8'b11010000;
    mem[97] <= 8'b11101111;
    mem[98] <= 8'b10101010;
    mem[99] <= 8'b11111011;
    mem[100] <= 8'b01000011;
    mem[101] <= 8'b01001101;
    mem[102] <= 8'b00110011;
    mem[103] <= 8'b10000101;
    mem[104] <= 8'b01000101;
    mem[105] <= 8'b11111001;
    mem[106] <= 8'b00000010;
    mem[107] <= 8'b01111111;
    mem[108] <= 8'b01010000;
    mem[109] <= 8'b00111100;
    mem[110] <= 8'b10011111;
    mem[111] <= 8'b10101000;
    mem[112] <= 8'b01010001;
    mem[113] <= 8'b10100011;
    mem[114] <= 8'b01000000;
    mem[115] <= 8'b10001111;
    mem[116] <= 8'b10010010;
    mem[117] <= 8'b10011101;
    mem[118] <= 8'b00111000;
    mem[119] <= 8'b11110101;
    mem[120] <= 8'b10111100;
    mem[121] <= 8'b10110110;
    mem[122] <= 8'b11011010;
    mem[123] <= 8'b00100001;
    mem[124] <= 8'b00010000;
    mem[125] <= 8'b11111111;
    mem[126] <= 8'b11110011;
    mem[127] <= 8'b11010010;
    mem[128] <= 8'b11001101;
    mem[129] <= 8'b00001100;
    mem[130] <= 8'b00010011;
    mem[131] <= 8'b11101100;
    mem[132] <= 8'b01011111;
    mem[133] <= 8'b10010111;
    mem[134] <= 8'b01000100;
    mem[135] <= 8'b00010111;
    mem[136] <= 8'b11000100;
    mem[137] <= 8'b10100111;
    mem[138] <= 8'b01111110;
    mem[139] <= 8'b00111101;
    mem[140] <= 8'b01100100;
    mem[141] <= 8'b01011101;
    mem[142] <= 8'b00011001;
    mem[143] <= 8'b01110011;
    mem[144] <= 8'b01100000;
    mem[145] <= 8'b10000001;
    mem[146] <= 8'b01001111;
    mem[147] <= 8'b11011100;
    mem[148] <= 8'b00100010;
    mem[149] <= 8'b00101010;
    mem[150] <= 8'b10010000;
    mem[151] <= 8'b10001000;
    mem[152] <= 8'b01000110;
    mem[153] <= 8'b11101110;
    mem[154] <= 8'b10111000;
    mem[155] <= 8'b00010100;
    mem[156] <= 8'b11011110;
    mem[157] <= 8'b01011110;
    mem[158] <= 8'b00001011;
    mem[159] <= 8'b11011011;
    mem[160] <= 8'b11100000;
    mem[161] <= 8'b00110010;
    mem[162] <= 8'b00111010;
    mem[163] <= 8'b00001010;
    mem[164] <= 8'b01001001;
    mem[165] <= 8'b00000110;
    mem[166] <= 8'b00100100;
    mem[167] <= 8'b01011100;
    mem[168] <= 8'b11000010;
    mem[169] <= 8'b11010011;
    mem[170] <= 8'b10101100;
    mem[171] <= 8'b01100010;
    mem[172] <= 8'b10010001;
    mem[173] <= 8'b10010101;
    mem[174] <= 8'b11100100;
    mem[175] <= 8'b01111001;
    mem[176] <= 8'b11100111;
    mem[177] <= 8'b11001000;
    mem[178] <= 8'b00110111;
    mem[179] <= 8'b01101101;
    mem[180] <= 8'b10001101;
    mem[181] <= 8'b11010101;
    mem[182] <= 8'b01001110;
    mem[183] <= 8'b10101001;
    mem[184] <= 8'b01101100;
    mem[185] <= 8'b01010110;
    mem[186] <= 8'b11110100;
    mem[187] <= 8'b11101010;
    mem[188] <= 8'b01100101;
    mem[189] <= 8'b01111010;
    mem[190] <= 8'b10101110;
    mem[191] <= 8'b00001000;
    mem[192] <= 8'b10111010;
    mem[193] <= 8'b01111000;
    mem[194] <= 8'b00100101;
    mem[195] <= 8'b00101110;
    mem[196] <= 8'b00011100;
    mem[197] <= 8'b10100110;
    mem[198] <= 8'b10110100;
    mem[199] <= 8'b11000110;
    mem[200] <= 8'b11101000;
    mem[201] <= 8'b11011101;
    mem[202] <= 8'b01110100;
    mem[203] <= 8'b00011111;
    mem[204] <= 8'b01001011;
    mem[205] <= 8'b10111101;
    mem[206] <= 8'b10001011;
    mem[207] <= 8'b10001010;
    mem[208] <= 8'b01110000;
    mem[209] <= 8'b00111110;
    mem[210] <= 8'b10110101;
    mem[211] <= 8'b01100110;
    mem[212] <= 8'b01001000;
    mem[213] <= 8'b00000011;
    mem[214] <= 8'b11110110;
    mem[215] <= 8'b00001110;
    mem[216] <= 8'b01100001;
    mem[217] <= 8'b00110101;
    mem[218] <= 8'b01010111;
    mem[219] <= 8'b10111001;
    mem[220] <= 8'b10000110;
    mem[221] <= 8'b11000001;
    mem[222] <= 8'b00011101;
    mem[223] <= 8'b10011110;
    mem[224] <= 8'b11100001;
    mem[225] <= 8'b11111000;
    mem[226] <= 8'b10011000;
    mem[227] <= 8'b00010001;
    mem[228] <= 8'b01101001;
    mem[229] <= 8'b11011001;
    mem[230] <= 8'b10001110;
    mem[231] <= 8'b10010100;
    mem[232] <= 8'b10011011;
    mem[233] <= 8'b00011110;
    mem[234] <= 8'b10000111;
    mem[235] <= 8'b11101001;
    mem[236] <= 8'b11001110;
    mem[237] <= 8'b01010101;
    mem[238] <= 8'b00101000;
    mem[239] <= 8'b11011111;
    mem[240] <= 8'b10001100;
    mem[241] <= 8'b10100001;
    mem[242] <= 8'b10001001;
    mem[243] <= 8'b00001101;
    mem[244] <= 8'b10111111;
    mem[245] <= 8'b11100110;
    mem[246] <= 8'b01000010;
    mem[247] <= 8'b01101000;
    mem[248] <= 8'b01000001;
    mem[249] <= 8'b10011001;
    mem[250] <= 8'b00101101;
    mem[251] <= 8'b00001111;
    mem[252] <= 8'b10110000;
    mem[253] <= 8'b01010100;
    mem[254] <= 8'b10111011;
    mem[255] <= 8'b00010110;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl_AES128_ENmgc_rom_19_512_8_1.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m112061603@ws34
//  Generated date: Sun Jun  9 02:20:57 2024
// ----------------------------------------------------------------------

// 
module AES128_ENmgc_rom_19_512_8_1 (addr, data_out, VDD, VSS
);
  input [8:0]addr ;
  output [7:0]data_out ;
  input VDD;
  input VSS;

  // Constants for ROM dimensions
  parameter n_width    = 8;
  parameter n_size     = 512;
  parameter n_numports = 1;
  parameter n_addr_w   = 9;
  parameter n_inreg    = 0;
  parameter n_outreg   = 0;

  // Declare storage for memory elements
  reg [7:0] mem [511:0];

  // Declare output registers
  reg [7:0] data_out_t;

  // Initialize ROM contents
  initial begin: rom_init_blk
    mem[0] <= 8'b00000000;
    mem[1] <= 8'b00000010;
    mem[2] <= 8'b00000100;
    mem[3] <= 8'b00000110;
    mem[4] <= 8'b00001000;
    mem[5] <= 8'b00001010;
    mem[6] <= 8'b00001100;
    mem[7] <= 8'b00001110;
    mem[8] <= 8'b00010000;
    mem[9] <= 8'b00010010;
    mem[10] <= 8'b00010100;
    mem[11] <= 8'b00010110;
    mem[12] <= 8'b00011000;
    mem[13] <= 8'b00011010;
    mem[14] <= 8'b00011100;
    mem[15] <= 8'b00011110;
    mem[16] <= 8'b00100000;
    mem[17] <= 8'b00100010;
    mem[18] <= 8'b00100100;
    mem[19] <= 8'b00100110;
    mem[20] <= 8'b00101000;
    mem[21] <= 8'b00101010;
    mem[22] <= 8'b00101100;
    mem[23] <= 8'b00101110;
    mem[24] <= 8'b00110000;
    mem[25] <= 8'b00110010;
    mem[26] <= 8'b00110100;
    mem[27] <= 8'b00110110;
    mem[28] <= 8'b00111000;
    mem[29] <= 8'b00111010;
    mem[30] <= 8'b00111100;
    mem[31] <= 8'b00111110;
    mem[32] <= 8'b01000000;
    mem[33] <= 8'b01000010;
    mem[34] <= 8'b01000100;
    mem[35] <= 8'b01000110;
    mem[36] <= 8'b01001000;
    mem[37] <= 8'b01001010;
    mem[38] <= 8'b01001100;
    mem[39] <= 8'b01001110;
    mem[40] <= 8'b01010000;
    mem[41] <= 8'b01010010;
    mem[42] <= 8'b01010100;
    mem[43] <= 8'b01010110;
    mem[44] <= 8'b01011000;
    mem[45] <= 8'b01011010;
    mem[46] <= 8'b01011100;
    mem[47] <= 8'b01011110;
    mem[48] <= 8'b01100000;
    mem[49] <= 8'b01100010;
    mem[50] <= 8'b01100100;
    mem[51] <= 8'b01100110;
    mem[52] <= 8'b01101000;
    mem[53] <= 8'b01101010;
    mem[54] <= 8'b01101100;
    mem[55] <= 8'b01101110;
    mem[56] <= 8'b01110000;
    mem[57] <= 8'b01110010;
    mem[58] <= 8'b01110100;
    mem[59] <= 8'b01110110;
    mem[60] <= 8'b01111000;
    mem[61] <= 8'b01111010;
    mem[62] <= 8'b01111100;
    mem[63] <= 8'b01111110;
    mem[64] <= 8'b10000000;
    mem[65] <= 8'b10000010;
    mem[66] <= 8'b10000100;
    mem[67] <= 8'b10000110;
    mem[68] <= 8'b10001000;
    mem[69] <= 8'b10001010;
    mem[70] <= 8'b10001100;
    mem[71] <= 8'b10001110;
    mem[72] <= 8'b10010000;
    mem[73] <= 8'b10010010;
    mem[74] <= 8'b10010100;
    mem[75] <= 8'b10010110;
    mem[76] <= 8'b10011000;
    mem[77] <= 8'b10011010;
    mem[78] <= 8'b10011100;
    mem[79] <= 8'b10011110;
    mem[80] <= 8'b10100000;
    mem[81] <= 8'b10100010;
    mem[82] <= 8'b10100100;
    mem[83] <= 8'b10100110;
    mem[84] <= 8'b10101000;
    mem[85] <= 8'b10101010;
    mem[86] <= 8'b10101100;
    mem[87] <= 8'b10101110;
    mem[88] <= 8'b10110000;
    mem[89] <= 8'b10110010;
    mem[90] <= 8'b10110100;
    mem[91] <= 8'b10110110;
    mem[92] <= 8'b10111000;
    mem[93] <= 8'b10111010;
    mem[94] <= 8'b10111100;
    mem[95] <= 8'b10111110;
    mem[96] <= 8'b11000000;
    mem[97] <= 8'b11000010;
    mem[98] <= 8'b11000100;
    mem[99] <= 8'b11000110;
    mem[100] <= 8'b11001000;
    mem[101] <= 8'b11001010;
    mem[102] <= 8'b11001100;
    mem[103] <= 8'b11001110;
    mem[104] <= 8'b11010000;
    mem[105] <= 8'b11010010;
    mem[106] <= 8'b11010100;
    mem[107] <= 8'b11010110;
    mem[108] <= 8'b11011000;
    mem[109] <= 8'b11011010;
    mem[110] <= 8'b11011100;
    mem[111] <= 8'b11011110;
    mem[112] <= 8'b11100000;
    mem[113] <= 8'b11100010;
    mem[114] <= 8'b11100100;
    mem[115] <= 8'b11100110;
    mem[116] <= 8'b11101000;
    mem[117] <= 8'b11101010;
    mem[118] <= 8'b11101100;
    mem[119] <= 8'b11101110;
    mem[120] <= 8'b11110000;
    mem[121] <= 8'b11110010;
    mem[122] <= 8'b11110100;
    mem[123] <= 8'b11110110;
    mem[124] <= 8'b11111000;
    mem[125] <= 8'b11111010;
    mem[126] <= 8'b11111100;
    mem[127] <= 8'b11111110;
    mem[128] <= 8'b00011011;
    mem[129] <= 8'b00011001;
    mem[130] <= 8'b00011111;
    mem[131] <= 8'b00011101;
    mem[132] <= 8'b00010011;
    mem[133] <= 8'b00010001;
    mem[134] <= 8'b00010111;
    mem[135] <= 8'b00010101;
    mem[136] <= 8'b00001011;
    mem[137] <= 8'b00001001;
    mem[138] <= 8'b00001111;
    mem[139] <= 8'b00001101;
    mem[140] <= 8'b00000011;
    mem[141] <= 8'b00000001;
    mem[142] <= 8'b00000111;
    mem[143] <= 8'b00000101;
    mem[144] <= 8'b00111011;
    mem[145] <= 8'b00111001;
    mem[146] <= 8'b00111111;
    mem[147] <= 8'b00111101;
    mem[148] <= 8'b00110011;
    mem[149] <= 8'b00110001;
    mem[150] <= 8'b00110111;
    mem[151] <= 8'b00110101;
    mem[152] <= 8'b00101011;
    mem[153] <= 8'b00101001;
    mem[154] <= 8'b00101111;
    mem[155] <= 8'b00101101;
    mem[156] <= 8'b00100011;
    mem[157] <= 8'b00100001;
    mem[158] <= 8'b00100111;
    mem[159] <= 8'b00100101;
    mem[160] <= 8'b01011011;
    mem[161] <= 8'b01011001;
    mem[162] <= 8'b01011111;
    mem[163] <= 8'b01011101;
    mem[164] <= 8'b01010011;
    mem[165] <= 8'b01010001;
    mem[166] <= 8'b01010111;
    mem[167] <= 8'b01010101;
    mem[168] <= 8'b01001011;
    mem[169] <= 8'b01001001;
    mem[170] <= 8'b01001111;
    mem[171] <= 8'b01001101;
    mem[172] <= 8'b01000011;
    mem[173] <= 8'b01000001;
    mem[174] <= 8'b01000111;
    mem[175] <= 8'b01000101;
    mem[176] <= 8'b01111011;
    mem[177] <= 8'b01111001;
    mem[178] <= 8'b01111111;
    mem[179] <= 8'b01111101;
    mem[180] <= 8'b01110011;
    mem[181] <= 8'b01110001;
    mem[182] <= 8'b01110111;
    mem[183] <= 8'b01110101;
    mem[184] <= 8'b01101011;
    mem[185] <= 8'b01101001;
    mem[186] <= 8'b01101111;
    mem[187] <= 8'b01101101;
    mem[188] <= 8'b01100011;
    mem[189] <= 8'b01100001;
    mem[190] <= 8'b01100111;
    mem[191] <= 8'b01100101;
    mem[192] <= 8'b10011011;
    mem[193] <= 8'b10011001;
    mem[194] <= 8'b10011111;
    mem[195] <= 8'b10011101;
    mem[196] <= 8'b10010011;
    mem[197] <= 8'b10010001;
    mem[198] <= 8'b10010111;
    mem[199] <= 8'b10010101;
    mem[200] <= 8'b10001011;
    mem[201] <= 8'b10001001;
    mem[202] <= 8'b10001111;
    mem[203] <= 8'b10001101;
    mem[204] <= 8'b10000011;
    mem[205] <= 8'b10000001;
    mem[206] <= 8'b10000111;
    mem[207] <= 8'b10000101;
    mem[208] <= 8'b10111011;
    mem[209] <= 8'b10111001;
    mem[210] <= 8'b10111111;
    mem[211] <= 8'b10111101;
    mem[212] <= 8'b10110011;
    mem[213] <= 8'b10110001;
    mem[214] <= 8'b10110111;
    mem[215] <= 8'b10110101;
    mem[216] <= 8'b10101011;
    mem[217] <= 8'b10101001;
    mem[218] <= 8'b10101111;
    mem[219] <= 8'b10101101;
    mem[220] <= 8'b10100011;
    mem[221] <= 8'b10100001;
    mem[222] <= 8'b10100111;
    mem[223] <= 8'b10100101;
    mem[224] <= 8'b11011011;
    mem[225] <= 8'b11011001;
    mem[226] <= 8'b11011111;
    mem[227] <= 8'b11011101;
    mem[228] <= 8'b11010011;
    mem[229] <= 8'b11010001;
    mem[230] <= 8'b11010111;
    mem[231] <= 8'b11010101;
    mem[232] <= 8'b11001011;
    mem[233] <= 8'b11001001;
    mem[234] <= 8'b11001111;
    mem[235] <= 8'b11001101;
    mem[236] <= 8'b11000011;
    mem[237] <= 8'b11000001;
    mem[238] <= 8'b11000111;
    mem[239] <= 8'b11000101;
    mem[240] <= 8'b11111011;
    mem[241] <= 8'b11111001;
    mem[242] <= 8'b11111111;
    mem[243] <= 8'b11111101;
    mem[244] <= 8'b11110011;
    mem[245] <= 8'b11110001;
    mem[246] <= 8'b11110111;
    mem[247] <= 8'b11110101;
    mem[248] <= 8'b11101011;
    mem[249] <= 8'b11101001;
    mem[250] <= 8'b11101111;
    mem[251] <= 8'b11101101;
    mem[252] <= 8'b11100011;
    mem[253] <= 8'b11100001;
    mem[254] <= 8'b11100111;
    mem[255] <= 8'b11100101;
    mem[256] <= 8'b00000000;
    mem[257] <= 8'b00000011;
    mem[258] <= 8'b00000110;
    mem[259] <= 8'b00000101;
    mem[260] <= 8'b00001100;
    mem[261] <= 8'b00001111;
    mem[262] <= 8'b00001010;
    mem[263] <= 8'b00001001;
    mem[264] <= 8'b00011000;
    mem[265] <= 8'b00011011;
    mem[266] <= 8'b00011110;
    mem[267] <= 8'b00011101;
    mem[268] <= 8'b00010100;
    mem[269] <= 8'b00010111;
    mem[270] <= 8'b00010010;
    mem[271] <= 8'b00010001;
    mem[272] <= 8'b00110000;
    mem[273] <= 8'b00110011;
    mem[274] <= 8'b00110110;
    mem[275] <= 8'b00110101;
    mem[276] <= 8'b00111100;
    mem[277] <= 8'b00111111;
    mem[278] <= 8'b00111010;
    mem[279] <= 8'b00111001;
    mem[280] <= 8'b00101000;
    mem[281] <= 8'b00101011;
    mem[282] <= 8'b00101110;
    mem[283] <= 8'b00101101;
    mem[284] <= 8'b00100100;
    mem[285] <= 8'b00100111;
    mem[286] <= 8'b00100010;
    mem[287] <= 8'b00100001;
    mem[288] <= 8'b01100000;
    mem[289] <= 8'b01100011;
    mem[290] <= 8'b01100110;
    mem[291] <= 8'b01100101;
    mem[292] <= 8'b01101100;
    mem[293] <= 8'b01101111;
    mem[294] <= 8'b01101010;
    mem[295] <= 8'b01101001;
    mem[296] <= 8'b01111000;
    mem[297] <= 8'b01111011;
    mem[298] <= 8'b01111110;
    mem[299] <= 8'b01111101;
    mem[300] <= 8'b01110100;
    mem[301] <= 8'b01110111;
    mem[302] <= 8'b01110010;
    mem[303] <= 8'b01110001;
    mem[304] <= 8'b01010000;
    mem[305] <= 8'b01010011;
    mem[306] <= 8'b01010110;
    mem[307] <= 8'b01010101;
    mem[308] <= 8'b01011100;
    mem[309] <= 8'b01011111;
    mem[310] <= 8'b01011010;
    mem[311] <= 8'b01011001;
    mem[312] <= 8'b01001000;
    mem[313] <= 8'b01001011;
    mem[314] <= 8'b01001110;
    mem[315] <= 8'b01001101;
    mem[316] <= 8'b01000100;
    mem[317] <= 8'b01000111;
    mem[318] <= 8'b01000010;
    mem[319] <= 8'b01000001;
    mem[320] <= 8'b11000000;
    mem[321] <= 8'b11000011;
    mem[322] <= 8'b11000110;
    mem[323] <= 8'b11000101;
    mem[324] <= 8'b11001100;
    mem[325] <= 8'b11001111;
    mem[326] <= 8'b11001010;
    mem[327] <= 8'b11001001;
    mem[328] <= 8'b11011000;
    mem[329] <= 8'b11011011;
    mem[330] <= 8'b11011110;
    mem[331] <= 8'b11011101;
    mem[332] <= 8'b11010100;
    mem[333] <= 8'b11010111;
    mem[334] <= 8'b11010010;
    mem[335] <= 8'b11010001;
    mem[336] <= 8'b11110000;
    mem[337] <= 8'b11110011;
    mem[338] <= 8'b11110110;
    mem[339] <= 8'b11110101;
    mem[340] <= 8'b11111100;
    mem[341] <= 8'b11111111;
    mem[342] <= 8'b11111010;
    mem[343] <= 8'b11111001;
    mem[344] <= 8'b11101000;
    mem[345] <= 8'b11101011;
    mem[346] <= 8'b11101110;
    mem[347] <= 8'b11101101;
    mem[348] <= 8'b11100100;
    mem[349] <= 8'b11100111;
    mem[350] <= 8'b11100010;
    mem[351] <= 8'b11100001;
    mem[352] <= 8'b10100000;
    mem[353] <= 8'b10100011;
    mem[354] <= 8'b10100110;
    mem[355] <= 8'b10100101;
    mem[356] <= 8'b10101100;
    mem[357] <= 8'b10101111;
    mem[358] <= 8'b10101010;
    mem[359] <= 8'b10101001;
    mem[360] <= 8'b10111000;
    mem[361] <= 8'b10111011;
    mem[362] <= 8'b10111110;
    mem[363] <= 8'b10111101;
    mem[364] <= 8'b10110100;
    mem[365] <= 8'b10110111;
    mem[366] <= 8'b10110010;
    mem[367] <= 8'b10110001;
    mem[368] <= 8'b10010000;
    mem[369] <= 8'b10010011;
    mem[370] <= 8'b10010110;
    mem[371] <= 8'b10010101;
    mem[372] <= 8'b10011100;
    mem[373] <= 8'b10011111;
    mem[374] <= 8'b10011010;
    mem[375] <= 8'b10011001;
    mem[376] <= 8'b10001000;
    mem[377] <= 8'b10001011;
    mem[378] <= 8'b10001110;
    mem[379] <= 8'b10001101;
    mem[380] <= 8'b10000100;
    mem[381] <= 8'b10000111;
    mem[382] <= 8'b10000010;
    mem[383] <= 8'b10000001;
    mem[384] <= 8'b10011011;
    mem[385] <= 8'b10011000;
    mem[386] <= 8'b10011101;
    mem[387] <= 8'b10011110;
    mem[388] <= 8'b10010111;
    mem[389] <= 8'b10010100;
    mem[390] <= 8'b10010001;
    mem[391] <= 8'b10010010;
    mem[392] <= 8'b10000011;
    mem[393] <= 8'b10000000;
    mem[394] <= 8'b10000101;
    mem[395] <= 8'b10000110;
    mem[396] <= 8'b10001111;
    mem[397] <= 8'b10001100;
    mem[398] <= 8'b10001001;
    mem[399] <= 8'b10001010;
    mem[400] <= 8'b10101011;
    mem[401] <= 8'b10101000;
    mem[402] <= 8'b10101101;
    mem[403] <= 8'b10101110;
    mem[404] <= 8'b10100111;
    mem[405] <= 8'b10100100;
    mem[406] <= 8'b10100001;
    mem[407] <= 8'b10100010;
    mem[408] <= 8'b10110011;
    mem[409] <= 8'b10110000;
    mem[410] <= 8'b10110101;
    mem[411] <= 8'b10110110;
    mem[412] <= 8'b10111111;
    mem[413] <= 8'b10111100;
    mem[414] <= 8'b10111001;
    mem[415] <= 8'b10111010;
    mem[416] <= 8'b11111011;
    mem[417] <= 8'b11111000;
    mem[418] <= 8'b11111101;
    mem[419] <= 8'b11111110;
    mem[420] <= 8'b11110111;
    mem[421] <= 8'b11110100;
    mem[422] <= 8'b11110001;
    mem[423] <= 8'b11110010;
    mem[424] <= 8'b11100011;
    mem[425] <= 8'b11100000;
    mem[426] <= 8'b11100101;
    mem[427] <= 8'b11100110;
    mem[428] <= 8'b11101111;
    mem[429] <= 8'b11101100;
    mem[430] <= 8'b11101001;
    mem[431] <= 8'b11101010;
    mem[432] <= 8'b11001011;
    mem[433] <= 8'b11001000;
    mem[434] <= 8'b11001101;
    mem[435] <= 8'b11001110;
    mem[436] <= 8'b11000111;
    mem[437] <= 8'b11000100;
    mem[438] <= 8'b11000001;
    mem[439] <= 8'b11000010;
    mem[440] <= 8'b11010011;
    mem[441] <= 8'b11010000;
    mem[442] <= 8'b11010101;
    mem[443] <= 8'b11010110;
    mem[444] <= 8'b11011111;
    mem[445] <= 8'b11011100;
    mem[446] <= 8'b11011001;
    mem[447] <= 8'b11011010;
    mem[448] <= 8'b01011011;
    mem[449] <= 8'b01011000;
    mem[450] <= 8'b01011101;
    mem[451] <= 8'b01011110;
    mem[452] <= 8'b01010111;
    mem[453] <= 8'b01010100;
    mem[454] <= 8'b01010001;
    mem[455] <= 8'b01010010;
    mem[456] <= 8'b01000011;
    mem[457] <= 8'b01000000;
    mem[458] <= 8'b01000101;
    mem[459] <= 8'b01000110;
    mem[460] <= 8'b01001111;
    mem[461] <= 8'b01001100;
    mem[462] <= 8'b01001001;
    mem[463] <= 8'b01001010;
    mem[464] <= 8'b01101011;
    mem[465] <= 8'b01101000;
    mem[466] <= 8'b01101101;
    mem[467] <= 8'b01101110;
    mem[468] <= 8'b01100111;
    mem[469] <= 8'b01100100;
    mem[470] <= 8'b01100001;
    mem[471] <= 8'b01100010;
    mem[472] <= 8'b01110011;
    mem[473] <= 8'b01110000;
    mem[474] <= 8'b01110101;
    mem[475] <= 8'b01110110;
    mem[476] <= 8'b01111111;
    mem[477] <= 8'b01111100;
    mem[478] <= 8'b01111001;
    mem[479] <= 8'b01111010;
    mem[480] <= 8'b00111011;
    mem[481] <= 8'b00111000;
    mem[482] <= 8'b00111101;
    mem[483] <= 8'b00111110;
    mem[484] <= 8'b00110111;
    mem[485] <= 8'b00110100;
    mem[486] <= 8'b00110001;
    mem[487] <= 8'b00110010;
    mem[488] <= 8'b00100011;
    mem[489] <= 8'b00100000;
    mem[490] <= 8'b00100101;
    mem[491] <= 8'b00100110;
    mem[492] <= 8'b00101111;
    mem[493] <= 8'b00101100;
    mem[494] <= 8'b00101001;
    mem[495] <= 8'b00101010;
    mem[496] <= 8'b00001011;
    mem[497] <= 8'b00001000;
    mem[498] <= 8'b00001101;
    mem[499] <= 8'b00001110;
    mem[500] <= 8'b00000111;
    mem[501] <= 8'b00000100;
    mem[502] <= 8'b00000001;
    mem[503] <= 8'b00000010;
    mem[504] <= 8'b00010011;
    mem[505] <= 8'b00010000;
    mem[506] <= 8'b00010101;
    mem[507] <= 8'b00010110;
    mem[508] <= 8'b00011111;
    mem[509] <= 8'b00011100;
    mem[510] <= 8'b00011001;
    mem[511] <= 8'b00011010;
  end


  // Combinational ROM read block
  always@(*)
  begin
    data_out_t <= mem[addr];
  end

  // Output register assignment
  assign data_out = data_out_t;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   m112061603@ws34
//  Generated date: Sun Jun  9 02:20:57 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module AES128_EN_run_run_fsm (
  clk, rst, arst_n, run_wen, fsm_output, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input run_wen;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input VDD;
  input VSS;

  // FSM State Type Declaration for AES128_EN_run_run_fsm_1
  parameter
    run_rlp_C_0 = 3'd0,
    main_C_0 = 3'd1,
    main_C_1 = 3'd2,
    main_C_2 = 3'd3,
    main_C_3 = 3'd4,
    main_C_4 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : AES128_EN_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 6'b000010;
        state_var_NS = main_C_1;
      end
      main_C_1 : begin
        fsm_output = 6'b000100;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 6'b001000;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 6'b010000;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 6'b100000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 6'b000001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( rst ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_staller
// ------------------------------------------------------------------


module AES128_EN_run_staller (
  clk, rst, arst_n, run_wen, plaintext_in_rsci_iden, plaintext_in_rsci_wen_comp,
      key_in_rsci_iden, key_in_rsci_wen_comp, ciphertext_out_rsci_iden, ciphertext_out_rsci_wen_comp,
      run_flen_unreg, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  output run_wen;
  input plaintext_in_rsci_iden;
  input plaintext_in_rsci_wen_comp;
  input key_in_rsci_iden;
  input key_in_rsci_wen_comp;
  input ciphertext_out_rsci_iden;
  input ciphertext_out_rsci_wen_comp;
  input run_flen_unreg;
  input VDD;
  input VSS;

  // Interconnect Declarations
  reg run_flen_shf_4;
  reg run_flen_shf_3;
  reg run_flen_shf_2;
  reg run_flen_shf_1;
  reg run_flen_shf_0;


  // Interconnect Declarations for Component Instantiations 
  assign run_wen = plaintext_in_rsci_wen_comp & key_in_rsci_wen_comp & ciphertext_out_rsci_wen_comp
      & (~(run_flen_shf_4 & run_flen_shf_3 & run_flen_shf_2 & run_flen_shf_1 & run_flen_shf_0
      & run_flen_unreg));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      run_flen_shf_4 <= 1'b0;
      run_flen_shf_3 <= 1'b0;
      run_flen_shf_2 <= 1'b0;
      run_flen_shf_1 <= 1'b0;
      run_flen_shf_0 <= 1'b0;
    end
    else if ( rst ) begin
      run_flen_shf_4 <= 1'b0;
      run_flen_shf_3 <= 1'b0;
      run_flen_shf_2 <= 1'b0;
      run_flen_shf_1 <= 1'b0;
      run_flen_shf_0 <= 1'b0;
    end
    else begin
      run_flen_shf_4 <= run_flen_shf_3;
      run_flen_shf_3 <= run_flen_shf_2;
      run_flen_shf_2 <= run_flen_shf_1;
      run_flen_shf_1 <= run_flen_shf_0;
      run_flen_shf_0 <= run_flen_unreg & (~(plaintext_in_rsci_iden | key_in_rsci_iden
          | ciphertext_out_rsci_iden));
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_dp
// ------------------------------------------------------------------


module AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_dp (
  clk, rst, arst_n, ciphertext_out_rsci_oswt_unreg, ciphertext_out_rsci_bawt, ciphertext_out_rsci_iden,
      ciphertext_out_rsci_wen_comp, ciphertext_out_rsci_biwt, ciphertext_out_rsci_bdwt,
      ciphertext_out_rsci_bcwt, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input ciphertext_out_rsci_oswt_unreg;
  output ciphertext_out_rsci_bawt;
  output ciphertext_out_rsci_iden;
  output ciphertext_out_rsci_wen_comp;
  input ciphertext_out_rsci_biwt;
  input ciphertext_out_rsci_bdwt;
  output ciphertext_out_rsci_bcwt;
  reg ciphertext_out_rsci_bcwt;
  input VDD;
  input VSS;


  // Interconnect Declarations for Component Instantiations 
  assign ciphertext_out_rsci_iden = ciphertext_out_rsci_biwt | ciphertext_out_rsci_bdwt;
  assign ciphertext_out_rsci_bawt = ciphertext_out_rsci_biwt | ciphertext_out_rsci_bcwt;
  assign ciphertext_out_rsci_wen_comp = (~ ciphertext_out_rsci_oswt_unreg) | ciphertext_out_rsci_bawt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ciphertext_out_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      ciphertext_out_rsci_bcwt <= 1'b0;
    end
    else begin
      ciphertext_out_rsci_bcwt <= ~((~(ciphertext_out_rsci_bcwt | ciphertext_out_rsci_biwt))
          | ciphertext_out_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_ctrl
// ------------------------------------------------------------------


module AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_ctrl (
  run_wen, ciphertext_out_rsci_oswt_unreg, ciphertext_out_rsci_iswt0, ciphertext_out_rsci_biwt,
      ciphertext_out_rsci_bdwt, ciphertext_out_rsci_bcwt, ciphertext_out_rsci_irdy,
      ciphertext_out_rsci_ivld_run_sct, VDD, VSS
);
  input run_wen;
  input ciphertext_out_rsci_oswt_unreg;
  input ciphertext_out_rsci_iswt0;
  output ciphertext_out_rsci_biwt;
  output ciphertext_out_rsci_bdwt;
  input ciphertext_out_rsci_bcwt;
  input ciphertext_out_rsci_irdy;
  output ciphertext_out_rsci_ivld_run_sct;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire ciphertext_out_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ciphertext_out_rsci_bdwt = ciphertext_out_rsci_oswt_unreg & run_wen;
  assign ciphertext_out_rsci_biwt = ciphertext_out_rsci_ogwt & ciphertext_out_rsci_irdy;
  assign ciphertext_out_rsci_ogwt = ciphertext_out_rsci_iswt0 & (~ ciphertext_out_rsci_bcwt);
  assign ciphertext_out_rsci_ivld_run_sct = ciphertext_out_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_key_in_rsci_key_in_wait_dp
// ------------------------------------------------------------------


module AES128_EN_run_key_in_rsci_key_in_wait_dp (
  clk, rst, arst_n, key_in_rsci_oswt_unreg, key_in_rsci_bawt, key_in_rsci_iden, key_in_rsci_wen_comp,
      key_in_rsci_idat_mxwt, key_in_rsci_biwt, key_in_rsci_bdwt, key_in_rsci_bcwt,
      key_in_rsci_idat, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input key_in_rsci_oswt_unreg;
  output key_in_rsci_bawt;
  output key_in_rsci_iden;
  output key_in_rsci_wen_comp;
  output [127:0] key_in_rsci_idat_mxwt;
  input key_in_rsci_biwt;
  input key_in_rsci_bdwt;
  output key_in_rsci_bcwt;
  reg key_in_rsci_bcwt;
  input [127:0] key_in_rsci_idat;
  input VDD;
  input VSS;

  // Interconnect Declarations
  reg [127:0] key_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign key_in_rsci_iden = key_in_rsci_biwt | key_in_rsci_bdwt;
  assign key_in_rsci_bawt = key_in_rsci_biwt | key_in_rsci_bcwt;
  assign key_in_rsci_wen_comp = (~ key_in_rsci_oswt_unreg) | key_in_rsci_bawt;
  assign key_in_rsci_idat_mxwt = MUX_v_128_2_2(key_in_rsci_idat, key_in_rsci_idat_bfwt,
      key_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      key_in_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      key_in_rsci_bcwt <= 1'b0;
    end
    else begin
      key_in_rsci_bcwt <= ~((~(key_in_rsci_bcwt | key_in_rsci_biwt)) | key_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( key_in_rsci_biwt ) begin
      key_in_rsci_idat_bfwt <= key_in_rsci_idat;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_key_in_rsci_key_in_wait_ctrl
// ------------------------------------------------------------------


module AES128_EN_run_key_in_rsci_key_in_wait_ctrl (
  run_wen, key_in_rsci_oswt_unreg, key_in_rsci_iswt0, key_in_rsci_biwt, key_in_rsci_bdwt,
      key_in_rsci_bcwt, key_in_rsci_irdy_run_sct, key_in_rsci_ivld, VDD, VSS
);
  input run_wen;
  input key_in_rsci_oswt_unreg;
  input key_in_rsci_iswt0;
  output key_in_rsci_biwt;
  output key_in_rsci_bdwt;
  input key_in_rsci_bcwt;
  output key_in_rsci_irdy_run_sct;
  input key_in_rsci_ivld;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire key_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign key_in_rsci_bdwt = key_in_rsci_oswt_unreg & run_wen;
  assign key_in_rsci_biwt = key_in_rsci_ogwt & key_in_rsci_ivld;
  assign key_in_rsci_ogwt = key_in_rsci_iswt0 & (~ key_in_rsci_bcwt);
  assign key_in_rsci_irdy_run_sct = key_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_dp
// ------------------------------------------------------------------


module AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_dp (
  clk, rst, arst_n, plaintext_in_rsci_oswt_unreg, plaintext_in_rsci_bawt, plaintext_in_rsci_iden,
      plaintext_in_rsci_wen_comp, plaintext_in_rsci_idat_mxwt, plaintext_in_rsci_biwt,
      plaintext_in_rsci_bdwt, plaintext_in_rsci_bcwt, plaintext_in_rsci_idat, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input plaintext_in_rsci_oswt_unreg;
  output plaintext_in_rsci_bawt;
  output plaintext_in_rsci_iden;
  output plaintext_in_rsci_wen_comp;
  output [127:0] plaintext_in_rsci_idat_mxwt;
  input plaintext_in_rsci_biwt;
  input plaintext_in_rsci_bdwt;
  output plaintext_in_rsci_bcwt;
  reg plaintext_in_rsci_bcwt;
  input [127:0] plaintext_in_rsci_idat;
  input VDD;
  input VSS;

  // Interconnect Declarations
  reg [127:0] plaintext_in_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign plaintext_in_rsci_iden = plaintext_in_rsci_biwt | plaintext_in_rsci_bdwt;
  assign plaintext_in_rsci_bawt = plaintext_in_rsci_biwt | plaintext_in_rsci_bcwt;
  assign plaintext_in_rsci_wen_comp = (~ plaintext_in_rsci_oswt_unreg) | plaintext_in_rsci_bawt;
  assign plaintext_in_rsci_idat_mxwt = MUX_v_128_2_2(plaintext_in_rsci_idat, plaintext_in_rsci_idat_bfwt,
      plaintext_in_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      plaintext_in_rsci_bcwt <= 1'b0;
    end
    else if ( rst ) begin
      plaintext_in_rsci_bcwt <= 1'b0;
    end
    else begin
      plaintext_in_rsci_bcwt <= ~((~(plaintext_in_rsci_bcwt | plaintext_in_rsci_biwt))
          | plaintext_in_rsci_bdwt);
    end
  end
  always @(posedge clk) begin
    if ( plaintext_in_rsci_biwt ) begin
      plaintext_in_rsci_idat_bfwt <= plaintext_in_rsci_idat;
    end
  end

  function automatic [127:0] MUX_v_128_2_2;
    input [127:0] input_0;
    input [127:0] input_1;
    input  sel;
    reg [127:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_128_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_ctrl
// ------------------------------------------------------------------


module AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_ctrl (
  run_wen, plaintext_in_rsci_oswt_unreg, plaintext_in_rsci_iswt0, plaintext_in_rsci_biwt,
      plaintext_in_rsci_bdwt, plaintext_in_rsci_bcwt, plaintext_in_rsci_irdy_run_sct,
      plaintext_in_rsci_ivld, VDD, VSS
);
  input run_wen;
  input plaintext_in_rsci_oswt_unreg;
  input plaintext_in_rsci_iswt0;
  output plaintext_in_rsci_biwt;
  output plaintext_in_rsci_bdwt;
  input plaintext_in_rsci_bcwt;
  output plaintext_in_rsci_irdy_run_sct;
  input plaintext_in_rsci_ivld;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire plaintext_in_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign plaintext_in_rsci_bdwt = plaintext_in_rsci_oswt_unreg & run_wen;
  assign plaintext_in_rsci_biwt = plaintext_in_rsci_ogwt & plaintext_in_rsci_ivld;
  assign plaintext_in_rsci_ogwt = plaintext_in_rsci_iswt0 & (~ plaintext_in_rsci_bcwt);
  assign plaintext_in_rsci_irdy_run_sct = plaintext_in_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_ciphertext_out_rsci
// ------------------------------------------------------------------


module AES128_EN_run_ciphertext_out_rsci (
  clk, rst, arst_n, ciphertext_out_rsc_dat, ciphertext_out_rsc_vld, ciphertext_out_rsc_rdy,
      run_wen, ciphertext_out_rsci_oswt_unreg, ciphertext_out_rsci_bawt, ciphertext_out_rsci_iden,
      ciphertext_out_rsci_iswt0, ciphertext_out_rsci_wen_comp, ciphertext_out_rsci_idat, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  output [127:0] ciphertext_out_rsc_dat;
  output ciphertext_out_rsc_vld;
  input ciphertext_out_rsc_rdy;
  input run_wen;
  input ciphertext_out_rsci_oswt_unreg;
  output ciphertext_out_rsci_bawt;
  output ciphertext_out_rsci_iden;
  input ciphertext_out_rsci_iswt0;
  output ciphertext_out_rsci_wen_comp;
  input [127:0] ciphertext_out_rsci_idat;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire ciphertext_out_rsci_biwt;
  wire ciphertext_out_rsci_bdwt;
  wire ciphertext_out_rsci_bcwt;
  wire ciphertext_out_rsci_irdy;
  wire ciphertext_out_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd128)) ciphertext_out_rsci (
      .irdy(ciphertext_out_rsci_irdy),
      .ivld(ciphertext_out_rsci_ivld_run_sct),
      .idat(ciphertext_out_rsci_idat),
      .rdy(ciphertext_out_rsc_rdy),
      .vld(ciphertext_out_rsc_vld),
      .dat(ciphertext_out_rsc_dat),
      .VDD(VDD),
      .VSS(VSS)
    );
  AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_ctrl AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .ciphertext_out_rsci_oswt_unreg(ciphertext_out_rsci_oswt_unreg),
      .ciphertext_out_rsci_iswt0(ciphertext_out_rsci_iswt0),
      .ciphertext_out_rsci_biwt(ciphertext_out_rsci_biwt),
      .ciphertext_out_rsci_bdwt(ciphertext_out_rsci_bdwt),
      .ciphertext_out_rsci_bcwt(ciphertext_out_rsci_bcwt),
      .ciphertext_out_rsci_irdy(ciphertext_out_rsci_irdy),
      .ciphertext_out_rsci_ivld_run_sct(ciphertext_out_rsci_ivld_run_sct),
      .VDD(VDD),
      .VSS(VSS)
    );
  AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_dp AES128_EN_run_ciphertext_out_rsci_ciphertext_out_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ciphertext_out_rsci_oswt_unreg(ciphertext_out_rsci_oswt_unreg),
      .ciphertext_out_rsci_bawt(ciphertext_out_rsci_bawt),
      .ciphertext_out_rsci_iden(ciphertext_out_rsci_iden),
      .ciphertext_out_rsci_wen_comp(ciphertext_out_rsci_wen_comp),
      .ciphertext_out_rsci_biwt(ciphertext_out_rsci_biwt),
      .ciphertext_out_rsci_bdwt(ciphertext_out_rsci_bdwt),
      .ciphertext_out_rsci_bcwt(ciphertext_out_rsci_bcwt),
      .VDD(VDD),
      .VSS(VSS)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_key_in_rsci
// ------------------------------------------------------------------


module AES128_EN_run_key_in_rsci (
  clk, rst, arst_n, key_in_rsc_dat, key_in_rsc_vld, key_in_rsc_rdy, run_wen, key_in_rsci_oswt_unreg,
      key_in_rsci_bawt, key_in_rsci_iden, key_in_rsci_iswt0, key_in_rsci_wen_comp,
      key_in_rsci_idat_mxwt, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input [127:0] key_in_rsc_dat;
  input key_in_rsc_vld;
  output key_in_rsc_rdy;
  input run_wen;
  input key_in_rsci_oswt_unreg;
  output key_in_rsci_bawt;
  output key_in_rsci_iden;
  input key_in_rsci_iswt0;
  output key_in_rsci_wen_comp;
  output [127:0] key_in_rsci_idat_mxwt;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire key_in_rsci_biwt;
  wire key_in_rsci_bdwt;
  wire key_in_rsci_bcwt;
  wire key_in_rsci_irdy_run_sct;
  wire key_in_rsci_ivld;
  wire [127:0] key_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd128)) key_in_rsci (
      .rdy(key_in_rsc_rdy),
      .vld(key_in_rsc_vld),
      .dat(key_in_rsc_dat),
      .irdy(key_in_rsci_irdy_run_sct),
      .ivld(key_in_rsci_ivld),
      .idat(key_in_rsci_idat),
      .VDD(VDD),
      .VSS(VSS)
    );
  AES128_EN_run_key_in_rsci_key_in_wait_ctrl AES128_EN_run_key_in_rsci_key_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .key_in_rsci_oswt_unreg(key_in_rsci_oswt_unreg),
      .key_in_rsci_iswt0(key_in_rsci_iswt0),
      .key_in_rsci_biwt(key_in_rsci_biwt),
      .key_in_rsci_bdwt(key_in_rsci_bdwt),
      .key_in_rsci_bcwt(key_in_rsci_bcwt),
      .key_in_rsci_irdy_run_sct(key_in_rsci_irdy_run_sct),
      .key_in_rsci_ivld(key_in_rsci_ivld),
      .VDD(VDD),
      .VSS(VSS)
    );
  AES128_EN_run_key_in_rsci_key_in_wait_dp AES128_EN_run_key_in_rsci_key_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .key_in_rsci_oswt_unreg(key_in_rsci_oswt_unreg),
      .key_in_rsci_bawt(key_in_rsci_bawt),
      .key_in_rsci_iden(key_in_rsci_iden),
      .key_in_rsci_wen_comp(key_in_rsci_wen_comp),
      .key_in_rsci_idat_mxwt(key_in_rsci_idat_mxwt),
      .key_in_rsci_biwt(key_in_rsci_biwt),
      .key_in_rsci_bdwt(key_in_rsci_bdwt),
      .key_in_rsci_bcwt(key_in_rsci_bcwt),
      .key_in_rsci_idat(key_in_rsci_idat),
      .VDD(VDD),
      .VSS(VSS)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run_plaintext_in_rsci
// ------------------------------------------------------------------


module AES128_EN_run_plaintext_in_rsci (
  clk, rst, arst_n, plaintext_in_rsc_dat, plaintext_in_rsc_vld, plaintext_in_rsc_rdy,
      run_wen, plaintext_in_rsci_oswt_unreg, plaintext_in_rsci_bawt, plaintext_in_rsci_iden,
      plaintext_in_rsci_iswt0, plaintext_in_rsci_wen_comp, plaintext_in_rsci_idat_mxwt, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input [127:0] plaintext_in_rsc_dat;
  input plaintext_in_rsc_vld;
  output plaintext_in_rsc_rdy;
  input run_wen;
  input plaintext_in_rsci_oswt_unreg;
  output plaintext_in_rsci_bawt;
  output plaintext_in_rsci_iden;
  input plaintext_in_rsci_iswt0;
  output plaintext_in_rsci_wen_comp;
  output [127:0] plaintext_in_rsci_idat_mxwt;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire plaintext_in_rsci_biwt;
  wire plaintext_in_rsci_bdwt;
  wire plaintext_in_rsci_bcwt;
  wire plaintext_in_rsci_irdy_run_sct;
  wire plaintext_in_rsci_ivld;
  wire [127:0] plaintext_in_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd128)) plaintext_in_rsci (
      .rdy(plaintext_in_rsc_rdy),
      .vld(plaintext_in_rsc_vld),
      .dat(plaintext_in_rsc_dat),
      .irdy(plaintext_in_rsci_irdy_run_sct),
      .ivld(plaintext_in_rsci_ivld),
      .idat(plaintext_in_rsci_idat),
      .VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_ctrl AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .plaintext_in_rsci_oswt_unreg(plaintext_in_rsci_oswt_unreg),
      .plaintext_in_rsci_iswt0(plaintext_in_rsci_iswt0),
      .plaintext_in_rsci_biwt(plaintext_in_rsci_biwt),
      .plaintext_in_rsci_bdwt(plaintext_in_rsci_bdwt),
      .plaintext_in_rsci_bcwt(plaintext_in_rsci_bcwt),
      .plaintext_in_rsci_irdy_run_sct(plaintext_in_rsci_irdy_run_sct),
      .plaintext_in_rsci_ivld(plaintext_in_rsci_ivld),
      .VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_dp AES128_EN_run_plaintext_in_rsci_plaintext_in_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .plaintext_in_rsci_oswt_unreg(plaintext_in_rsci_oswt_unreg),
      .plaintext_in_rsci_bawt(plaintext_in_rsci_bawt),
      .plaintext_in_rsci_iden(plaintext_in_rsci_iden),
      .plaintext_in_rsci_wen_comp(plaintext_in_rsci_wen_comp),
      .plaintext_in_rsci_idat_mxwt(plaintext_in_rsci_idat_mxwt),
      .plaintext_in_rsci_biwt(plaintext_in_rsci_biwt),
      .plaintext_in_rsci_bdwt(plaintext_in_rsci_bdwt),
      .plaintext_in_rsci_bcwt(plaintext_in_rsci_bcwt),
      .plaintext_in_rsci_idat(plaintext_in_rsci_idat),
      .VDD(VDD),
.VSS(VSS)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN_run
// ------------------------------------------------------------------


module AES128_EN_run (
  clk, rst, arst_n, plaintext_in_rsc_dat, plaintext_in_rsc_vld, plaintext_in_rsc_rdy,
      key_in_rsc_dat, key_in_rsc_vld, key_in_rsc_rdy, ciphertext_out_rsc_dat, ciphertext_out_rsc_vld,
      ciphertext_out_rsc_rdy, VDD, VSS
);
  input clk;
  input rst;
  input arst_n;
  input [127:0] plaintext_in_rsc_dat;
  input plaintext_in_rsc_vld;
  output plaintext_in_rsc_rdy;
  input [127:0] key_in_rsc_dat;
  input key_in_rsc_vld;
  output key_in_rsc_rdy;
  output [127:0] ciphertext_out_rsc_dat;
  output ciphertext_out_rsc_vld;
  input ciphertext_out_rsc_rdy;
  input VDD;
  input VSS;

  // Interconnect Declarations
  wire run_wen;
  wire plaintext_in_rsci_bawt;
  wire plaintext_in_rsci_iden;
  wire plaintext_in_rsci_wen_comp;
  wire [127:0] plaintext_in_rsci_idat_mxwt;
  wire key_in_rsci_bawt;
  wire key_in_rsci_iden;
  wire key_in_rsci_wen_comp;
  wire [127:0] key_in_rsci_idat_mxwt;
  wire ciphertext_out_rsci_bawt;
  wire ciphertext_out_rsci_iden;
  reg ciphertext_out_rsci_iswt0;
  wire ciphertext_out_rsci_wen_comp;
  reg [7:0] ciphertext_out_rsci_idat_119_112;
  reg [7:0] ciphertext_out_rsci_idat_111_104;
  reg [7:0] ciphertext_out_rsci_idat_103_96;
  reg [1:0] ciphertext_out_rsci_idat_95_94;
  reg [1:0] ciphertext_out_rsci_idat_93_92;
  reg ciphertext_out_rsci_idat_91;
  reg [1:0] ciphertext_out_rsci_idat_90_89;
  reg ciphertext_out_rsci_idat_88;
  reg [7:0] ciphertext_out_rsci_idat_87_80;
  reg [7:0] ciphertext_out_rsci_idat_79_72;
  reg [7:0] ciphertext_out_rsci_idat_71_64;
  reg [1:0] ciphertext_out_rsci_idat_63_62;
  reg [1:0] ciphertext_out_rsci_idat_61_60;
  reg ciphertext_out_rsci_idat_59;
  reg [1:0] ciphertext_out_rsci_idat_58_57;
  reg ciphertext_out_rsci_idat_56;
  reg [7:0] ciphertext_out_rsci_idat_55_48;
  reg [7:0] ciphertext_out_rsci_idat_47_40;
  reg [7:0] ciphertext_out_rsci_idat_39_32;
  reg [1:0] ciphertext_out_rsci_idat_31_30;
  reg [1:0] ciphertext_out_rsci_idat_29_28;
  reg ciphertext_out_rsci_idat_27;
  reg [1:0] ciphertext_out_rsci_idat_26_25;
  reg ciphertext_out_rsci_idat_24;
  reg [7:0] ciphertext_out_rsci_idat_23_16;
  reg [7:0] ciphertext_out_rsci_idat_15_8;
  reg [7:0] ciphertext_out_rsci_idat_7_0;
  reg [1:0] ciphertext_out_rsci_idat_127_126;
  reg [1:0] ciphertext_out_rsci_idat_125_124;
  reg ciphertext_out_rsci_idat_123;
  reg [1:0] ciphertext_out_rsci_idat_122_121;
  reg ciphertext_out_rsci_idat_120;
  wire [5:0] fsm_output;
  wire ROUND_ROUND_and_tmp;
  wire or_dcpl;
  wire and_dcpl;
  wire or_tmp;
  wire or_tmp_19;
  wire and_dcpl_35;
  wire and_dcpl_36;
  wire or_dcpl_43;
  wire or_dcpl_45;
  wire or_dcpl_48;
  wire or_dcpl_49;
  wire and_dcpl_49;
  wire or_dcpl_66;
  wire or_dcpl_67;
  wire or_dcpl_76;
  wire or_dcpl_80;
  wire or_dcpl_83;
  wire or_dcpl_88;
  wire or_dcpl_90;
  wire or_dcpl_94;
  wire or_dcpl_110;
  wire or_tmp_49;
  wire or_tmp_55;
  wire or_tmp_98;
  wire or_tmp_99;
  wire or_tmp_103;
  wire or_tmp_107;
  wire or_tmp_111;
  wire or_tmp_115;
  wire or_tmp_118;
  wire or_tmp_145;
  wire and_110_cse;
  reg main_stage_v_4;
  reg main_stage_v_5;
  reg main_stage_v_3;
  reg main_stage_v_2;
  reg main_stage_v_1;
  reg main_stage_v;
  wire main_stage_v_5_mx1;
  reg ROUND_not_mdf_sva_st_1;
  reg exitL_exit_ROUND_sva;
  reg ROUND_not_mdf_sva_st;
  reg ROUND_asn_itm;
  wire and_546_cse;
  wire AES128_EN_GenRoundKey_for_and_cse;
  wire ROUND_r_and_cse;
  wire state_arr_and_2_cse;
  wire state_arr_and_4_cse;
  wire roundkeys_and_cse;
  wire AES128_EN_ShiftRows_a_arr_and_cse;
  wire AES128_EN_MixColumns_for_for_for_else_and_1_cse;
  wire AES128_EN_ShiftRows_a_arr_and_1_cse;
  wire AES128_EN_MixColumns_for_for_for_else_and_2_cse;
  wire AES128_EN_ShiftRows_a_arr_and_11_cse;
  wire ROUND_and_2_cse;
  wire AES128_EN_MixColumns_for_for_for_else_and_7_cse;
  wire ROUND_and_9_cse;
  wire AES128_EN_AddRoundKey_2_for_for_and_cse;
  wire AES128_EN_GenRoundKey_1_for_and_cse;
  wire state_arr_and_3_cse;
  wire AES128_EN_AddRoundKey_2_for_for_and_15_cse;
  wire or_cse;
  wire nor_17_cse;
  wire and_10_cse;
  wire nor_8_cse;
  wire nand_26_cse;
  reg reg_key_in_rsci_iswt0_cse;
  wire and_20_cse;
  wire [7:0] data_out_out;
  wire [7:0] data_out_out_1;
  wire [7:0] data_out_out_2;
  wire [7:0] data_out_out_3;
  wire [7:0] data_out_out_4;
  wire [7:0] data_out_out_5;
  wire [7:0] data_out_out_6;
  wire [7:0] data_out_out_7;
  wire [7:0] data_out_out_8;
  wire [7:0] data_out_out_9;
  wire [7:0] data_out_out_10;
  wire [7:0] data_out_out_11;
  wire [7:0] data_out_out_12;
  wire [7:0] data_out_out_13;
  wire [7:0] data_out_out_14;
  wire [7:0] data_out_out_15;
  wire [7:0] data_out_out_16;
  wire [7:0] data_out_out_17;
  wire [7:0] data_out_out_18;
  reg [7:0] roundkeys_12_lpi_1;
  reg [7:0] roundkeys_13_lpi_1;
  reg [7:0] roundkeys_14_lpi_1;
  reg [7:0] roundkeys_15_lpi_1;
  reg [7:0] state_arr_1_3_1_lpi_1;
  reg [7:0] state_arr_2_0_1_lpi_1;
  reg [7:0] state_arr_2_1_1_lpi_1;
  reg [7:0] state_arr_1_0_1_lpi_1;
  reg [7:0] state_arr_3_2_1_lpi_1;
  reg [7:0] state_arr_0_0_lpi_1;
  reg [7:0] state_arr_3_3_1_lpi_1;
  reg [7:0] AES128_EN_ShiftRows_a_arr_0_0_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_2_0_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_1_3_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_2_1_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_1_2_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_2_2_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_1_1_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_2_3_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_1_0_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_3_0_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_0_3_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_3_1_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_0_2_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_3_2_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_0_1_sva;
  reg [7:0] AES128_EN_ShiftRows_a_arr_3_3_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  reg [3:0] ROUND_r_3_0_sva_1;
  reg AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_3_sva;
  reg [1:0] AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_2_1_sva;
  reg [1:0] AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_5_4_sva;
  reg AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_0_sva;
  reg [1:0] AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_7_6_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_3_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
  reg [7:0] AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva;
  reg [7:0] ROUND_mux_itm;
  reg [7:0] ROUND_mux_29_itm;
  reg [7:0] ROUND_mux_30_itm;
  reg [7:0] ROUND_mux_26_itm;
  reg [7:0] ROUND_mux_25_itm;
  reg [7:0] ROUND_mux_24_itm;
  reg [7:0] ROUND_mux_34_itm;
  reg [7:0] ROUND_mux_31_itm;
  reg [7:0] ROUND_mux_20_itm;
  reg [7:0] AES128_EN_Rcon_mux_itm;
  reg [7:0] ROUND_mux_2_itm;
  reg [7:0] ROUND_mux_3_itm;
  reg [7:0] ROUND_mux_6_itm;
  reg [7:0] ROUND_mux_7_itm;
  reg [7:0] ROUND_mux_10_itm;
  reg [7:0] ROUND_mux_11_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_24_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_18_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_19_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_16_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_8_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_4_itm;
  reg [7:0] AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_5_itm;
  reg [7:0] AES128_EN_AddRoundKey_2_for_2_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [7:0] AES128_EN_AddRoundKey_2_for_4_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
  reg [7:0] AES128_EN_AddRoundKey_2_for_2_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
  reg [7:0] AES128_EN_AddRoundKey_2_for_2_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
  reg AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_7_6;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_5_4;
  reg AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_3;
  reg [1:0] AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_2_1;
  reg AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_0;
  wire [3:0] ROUND_r_3_0_sva_2;
  wire [4:0] nl_ROUND_r_3_0_sva_2;
  wire [7:0] AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1;
  wire [7:0] AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1;
  wire [7:0] state_arr_0_1_1_sva_2;
  wire [7:0] state_arr_3_1_1_sva_2;
  wire [7:0] state_arr_0_2_1_sva_2;
  wire [7:0] state_arr_3_0_1_sva_2;
  wire [7:0] state_arr_0_3_1_sva_2;
  wire [7:0] state_arr_1_1_1_sva_2;
  wire [7:0] state_arr_1_2_1_sva_2;
  wire [7:0] state_arr_2_3_1_sva_2;
  wire [7:0] state_arr_2_2_1_sva_2;
  wire [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0;
  wire [7:0] AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva_mx1w0;
  wire main_stage_v_5_mx0c0;
  wire [3:0] ROUND_r_3_0_lpi_1_dfm_mx0;
  wire [7:0] xor_cse;
  wire [7:0] xor_cse_13;
  wire [7:0] xor_cse_14;
  wire [7:0] xor_cse_15;
  wire [7:0] xor_cse_16;
  wire [7:0] xor_cse_22;
  wire xor_cse_27;
  wire [1:0] xor_cse_34;
  wire xor_cse_41;
  wire [1:0] xor_cse_48;
  wire [1:0] xor_cse_55;
  wire [7:0] xor_cse_69;
  wire [7:0] xor_cse_72;
  wire AES128_EN_MixColumns_for_for_for_else_nor_1_cse;
  wire AES128_EN_SubBytes_1_for_for_and_cse;
  wire AES128_EN_SubBytes_1_for_for_and_1_cse;
  wire AES128_EN_MixColumns_for_for_for_else_or_cse;
  wire AES128_EN_MixColumns_for_for_for_else_or_1_cse;

  wire AES128_EN_GenRoundKey_for_mux_33_nl;
  wire or_139_nl;
  wire roundkeys_mux_nl;
  wire or_145_nl;
  wire roundkeys_mux_3_nl;
  wire or_148_nl;
  wire AES128_EN_ShiftRows_a_arr_mux_27_nl;
  wire or_154_nl;
  wire or_156_nl;
  wire AES128_EN_MixColumns_for_for_for_else_mux_18_nl;
  wire or_134_nl;
  wire AES128_EN_ShiftRows_a_arr_mux_28_nl;
  wire or_162_nl;
  wire AES128_EN_ShiftRows_a_arr_mux_29_nl;
  wire or_164_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_1_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_4_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_4_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_2_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_2_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire ROUND_mux_53_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_2_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_3_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_3_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire[7:0] AES128_EN_AddRoundKey_for_1_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire AES128_EN_ShiftRows_a_arr_mux_31_nl;
  wire[7:0] for_1_mux_8_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_12_rg_addr;
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_12_rg_addr = MUX1HOT_v_8_3_2(state_arr_3_0_1_sva_2,
      state_arr_1_2_1_sva_2, state_arr_0_2_1_sva_2, {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[3])});
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_11_rg_addr;
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_11_rg_addr = MUX_v_8_2_2(state_arr_2_3_1_sva_2,
      state_arr_0_3_1_sva_2, fsm_output[3]);
  wire[7:0] AES128_EN_AddRoundKey_for_4_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_7_rg_addr;
  assign AES128_EN_AddRoundKey_for_4_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[71:64]) ^ (key_in_rsci_idat_mxwt[71:64]);
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_7_rg_addr = MUX1HOT_v_8_6_2(state_arr_2_0_1_lpi_1,
      state_arr_1_3_1_lpi_1, ROUND_mux_34_itm, AES128_EN_ShiftRows_a_arr_1_0_sva,
      AES128_EN_AddRoundKey_for_4_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl, roundkeys_15_lpi_1,
      {(fsm_output[5]) , (fsm_output[4]) , (fsm_output[2]) , AES128_EN_SubBytes_1_for_for_and_cse
      , AES128_EN_SubBytes_1_for_for_and_1_cse , (fsm_output[3])});
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_1_rg_addr;
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_1_rg_addr = MUX1HOT_v_8_3_2(state_arr_3_1_1_sva_2,
      state_arr_1_1_1_sva_2, state_arr_0_1_1_sva_2, {(fsm_output[5]) , (fsm_output[4])
      , (fsm_output[3])});
  wire[7:0] AES128_EN_AddRoundKey_for_3_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_15_rg_addr;
  assign AES128_EN_AddRoundKey_for_3_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[79:72]) ^ (key_in_rsci_idat_mxwt[79:72]);
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_15_rg_addr = MUX1HOT_v_8_5_2(state_arr_1_0_1_lpi_1,
      ROUND_mux_31_itm, state_arr_3_3_1_lpi_1, state_arr_2_1_1_lpi_1, AES128_EN_AddRoundKey_for_3_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl,
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , AES128_EN_SubBytes_1_for_for_and_cse
      , AES128_EN_SubBytes_1_for_for_and_1_cse});
  wire[7:0] AES128_EN_AddRoundKey_for_2_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_10_rg_addr;
  assign AES128_EN_AddRoundKey_for_2_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[119:112]) ^ (key_in_rsci_idat_mxwt[119:112]);
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_10_rg_addr = MUX1HOT_v_8_6_2(state_arr_2_2_1_sva_2,
      ROUND_mux_30_itm, state_arr_1_0_1_lpi_1, AES128_EN_AddRoundKey_for_2_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl,
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva_mx1w0,
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva, {(fsm_output[5])
      , (fsm_output[2]) , AES128_EN_SubBytes_1_for_for_and_cse , AES128_EN_SubBytes_1_for_for_and_1_cse
      , (fsm_output[3]) , (fsm_output[4])});
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_rg_addr;
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_rg_addr = MUX1HOT_v_8_5_2(state_arr_2_1_1_lpi_1,
      ROUND_mux_25_itm, state_arr_0_0_lpi_1, roundkeys_12_lpi_1, (key_in_rsci_idat_mxwt[31:24]),
      {(fsm_output[5]) , (fsm_output[2]) , (fsm_output[4]) , AES128_EN_SubBytes_1_for_for_and_cse
      , AES128_EN_SubBytes_1_for_for_and_1_cse});
  wire[7:0] AES128_EN_AddRoundKey_for_3_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_14_rg_addr;
  assign AES128_EN_AddRoundKey_for_3_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[111:104]) ^ (key_in_rsci_idat_mxwt[111:104]);
  assign nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_14_rg_addr = MUX1HOT_v_8_5_2(state_arr_3_2_1_lpi_1,
      state_arr_2_0_1_lpi_1, AES128_EN_AddRoundKey_for_3_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl,
      ROUND_mux_26_itm, AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_7_ncse_sva,
      {(fsm_output[5]) , AES128_EN_SubBytes_1_for_for_and_cse , AES128_EN_SubBytes_1_for_for_and_1_cse
      , (fsm_output[2]) , (fsm_output[4])});
  wire[7:0] AES128_EN_AddRoundKey_for_1_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_rg_addr;
  assign AES128_EN_AddRoundKey_for_1_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[63:56]) ^ (key_in_rsci_idat_mxwt[63:56]);
  assign nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_rg_addr = MUX1HOT_v_8_4_2(ROUND_mux_itm,
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_itm,
      AES128_EN_AddRoundKey_for_1_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl, roundkeys_13_lpi_1,
      {(fsm_output[2]) , AES128_EN_SubBytes_1_for_for_and_cse , AES128_EN_SubBytes_1_for_for_and_1_cse
      , (fsm_output[3])});
  wire[7:0] AES128_EN_AddRoundKey_for_4_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_10_rg_addr;
  assign AES128_EN_AddRoundKey_for_4_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[39:32]) ^ (key_in_rsci_idat_mxwt[39:32]);
  assign nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_10_rg_addr = MUX1HOT_v_8_5_2(ROUND_mux_29_itm,
      state_arr_3_2_1_lpi_1, AES128_EN_AddRoundKey_for_4_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl,
      roundkeys_14_lpi_1, AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva,
      {(fsm_output[2]) , AES128_EN_SubBytes_1_for_for_and_cse , AES128_EN_SubBytes_1_for_for_and_1_cse
      , (fsm_output[3]) , (fsm_output[4])});
  wire[7:0] AES128_EN_AddRoundKey_for_1_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl;
  wire [7:0] nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_1_rg_addr;
  assign AES128_EN_AddRoundKey_for_1_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[31:24]) ^ (key_in_rsci_idat_mxwt[31:24]);
  assign nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_1_rg_addr = MUX1HOT_v_8_4_2(ROUND_mux_24_itm,
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_16_itm,
      AES128_EN_AddRoundKey_for_1_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl, ROUND_mux_20_itm,
      {(fsm_output[2]) , AES128_EN_SubBytes_1_for_for_and_cse , AES128_EN_SubBytes_1_for_for_and_1_cse
      , (fsm_output[3])});
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_6_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_31_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_6_nl
      = (~((fsm_output[2]) | (fsm_output[5]))) | (fsm_output[1]) | (fsm_output[4]);
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_31_nl = MUX1HOT_v_8_3_2(data_out_out_10,
      data_out_out_8, AES128_EN_ShiftRows_a_arr_2_2_sva, {(fsm_output[1]) , (fsm_output[2])
      , AES128_EN_MixColumns_for_for_for_else_or_1_cse});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_6_nl
      , AES128_EN_MixColumns_for_for_for_else_mux1h_31_nl};
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_24_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_14_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_24_nl = MUX1HOT_v_8_3_2(data_out_out_9,
      AES128_EN_ShiftRows_a_arr_2_1_sva, AES128_EN_ShiftRows_a_arr_1_0_sva, {AES128_EN_MixColumns_for_for_for_else_or_cse
      , (fsm_output[4]) , (fsm_output[3])});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_14_rg_addr
      = {1'b0, AES128_EN_MixColumns_for_for_for_else_mux1h_24_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_5_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_32_nl;
  wire AES128_EN_MixColumns_for_for_for_else_or_3_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_5_nl
      = (~((fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]))) | (fsm_output[3:2]!=2'b00);
  assign AES128_EN_MixColumns_for_for_for_else_or_3_nl = (fsm_output[4:3]!=2'b00);
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_32_nl = MUX1HOT_v_8_3_2(data_out_out_2,
      AES128_EN_ShiftRows_a_arr_3_0_sva, AES128_EN_ShiftRows_a_arr_1_1_sva, {AES128_EN_MixColumns_for_for_for_else_or_cse
      , (fsm_output[5]) , AES128_EN_MixColumns_for_for_for_else_or_3_nl});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_5_nl
      , AES128_EN_MixColumns_for_for_for_else_mux1h_32_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_4_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_33_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_15_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_4_nl
      = AES128_EN_MixColumns_for_for_for_else_nor_1_cse | (fsm_output[4]) | (fsm_output[2]);
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_33_nl = MUX1HOT_v_8_3_2(AES128_EN_ShiftRows_a_arr_3_1_sva,
      AES128_EN_ShiftRows_a_arr_2_3_sva, AES128_EN_ShiftRows_a_arr_0_3_sva, {AES128_EN_MixColumns_for_for_for_else_or_1_cse
      , (fsm_output[2]) , (fsm_output[3])});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_15_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_4_nl
      , AES128_EN_MixColumns_for_for_for_else_mux1h_33_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_3_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_34_nl;
  wire AES128_EN_MixColumns_for_for_for_else_or_5_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_11_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_3_nl
      = (fsm_output[5:2]!=4'b0001);
  assign AES128_EN_MixColumns_for_for_for_else_or_5_nl = (fsm_output[3:2]!=2'b00);
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_34_nl = MUX1HOT_v_8_3_2(AES128_EN_ShiftRows_a_arr_2_0_sva,
      AES128_EN_ShiftRows_a_arr_1_3_sva, AES128_EN_ShiftRows_a_arr_3_3_sva, {(fsm_output[4])
      , AES128_EN_MixColumns_for_for_for_else_or_5_nl , (fsm_output[5])});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_11_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_3_nl
      , AES128_EN_MixColumns_for_for_for_else_mux1h_34_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_2_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_mux1h_35_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_23_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_2_nl
      = (fsm_output[5:1]!=5'b00100);
  assign AES128_EN_MixColumns_for_for_for_else_mux1h_35_nl = MUX1HOT_v_8_4_2(data_out_out_8,
      AES128_EN_ShiftRows_a_arr_0_1_sva, AES128_EN_ShiftRows_a_arr_2_1_sva, AES128_EN_ShiftRows_a_arr_0_2_sva,
      {AES128_EN_MixColumns_for_for_for_else_or_cse , (fsm_output[5]) , (fsm_output[4])
      , (fsm_output[3])});
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_23_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_2_nl
      , AES128_EN_MixColumns_for_for_for_else_mux1h_35_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_1_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_2_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_1_nl
      = AES128_EN_MixColumns_for_for_for_else_nor_1_cse | (fsm_output[2]);
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_2_nl
      = MUX_v_8_2_2(data_out_out_10, AES128_EN_ShiftRows_a_arr_2_3_sva, fsm_output[5]);
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_1_nl
      , AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_2_nl};
  wire AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_nl;
  wire[7:0] AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_3_nl;
  wire [8:0] nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_13_rg_addr;
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_nl
      = (fsm_output[5:3]!=3'b010);
  assign AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_3_nl
      = MUX_v_8_2_2(AES128_EN_ShiftRows_a_arr_1_2_sva, AES128_EN_ShiftRows_a_arr_3_2_sva,
      fsm_output[5]);
  assign nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_13_rg_addr
      = {AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_or_nl
      , AES128_EN_MixColumns_for_for_for_else_AES128_EN_MixColumns_for_for_for_else_mux_3_nl};
  wire [127:0] nl_AES128_EN_run_ciphertext_out_rsci_inst_ciphertext_out_rsci_idat;
  assign nl_AES128_EN_run_ciphertext_out_rsci_inst_ciphertext_out_rsci_idat = {ciphertext_out_rsci_idat_127_126
      , ciphertext_out_rsci_idat_125_124 , ciphertext_out_rsci_idat_123 , ciphertext_out_rsci_idat_122_121
      , ciphertext_out_rsci_idat_120 , ciphertext_out_rsci_idat_119_112 , ciphertext_out_rsci_idat_111_104
      , ciphertext_out_rsci_idat_103_96 , ciphertext_out_rsci_idat_95_94 , ciphertext_out_rsci_idat_93_92
      , ciphertext_out_rsci_idat_91 , ciphertext_out_rsci_idat_90_89 , ciphertext_out_rsci_idat_88
      , ciphertext_out_rsci_idat_87_80 , ciphertext_out_rsci_idat_79_72 , ciphertext_out_rsci_idat_71_64
      , ciphertext_out_rsci_idat_63_62 , ciphertext_out_rsci_idat_61_60 , ciphertext_out_rsci_idat_59
      , ciphertext_out_rsci_idat_58_57 , ciphertext_out_rsci_idat_56 , ciphertext_out_rsci_idat_55_48
      , ciphertext_out_rsci_idat_47_40 , ciphertext_out_rsci_idat_39_32 , ciphertext_out_rsci_idat_31_30
      , ciphertext_out_rsci_idat_29_28 , ciphertext_out_rsci_idat_27 , ciphertext_out_rsci_idat_26_25
      , ciphertext_out_rsci_idat_24 , ciphertext_out_rsci_idat_23_16 , ciphertext_out_rsci_idat_15_8
      , ciphertext_out_rsci_idat_7_0};
  wire nor_1_nl;
  wire nor_3_nl;
  wire nand_33_nl;
  wire nand_34_nl;
  wire nand_35_nl;
  wire or_179_nl;
  wire  nl_AES128_EN_run_staller_inst_run_flen_unreg;
  assign nor_1_nl = ~((~((main_stage_v & (~ (fsm_output[0]))) | (main_stage_v_1 &
      (~ (fsm_output[0]))) | (main_stage_v_2 & (~ (fsm_output[0]))) | (main_stage_v_3
      & (~ (fsm_output[0]))) | (main_stage_v_4 & ((~((fsm_output[0]) | (fsm_output[5])))
      | (or_dcpl_67 & (fsm_output[5])))))) | and_10_cse);
  assign nor_3_nl = ~((main_stage_v & (~(main_stage_v_1 | main_stage_v_2 | main_stage_v_3
      | main_stage_v_4 | main_stage_v_5_mx1)) & (plaintext_in_rsci_bawt | (~ ROUND_asn_itm))
      & (key_in_rsci_bawt | (~ ROUND_asn_itm)) & (ciphertext_out_rsci_bawt | (~(ROUND_not_mdf_sva_st_1
      & main_stage_v_5_mx1)))) | (main_stage_v_5 & or_cse));
  assign nand_33_nl = ~(main_stage_v_1 & (~(main_stage_v_2 | main_stage_v_3 | main_stage_v_4
      | main_stage_v_5)));
  assign nand_34_nl = ~(main_stage_v_2 & (~(main_stage_v_3 | main_stage_v_4 | main_stage_v_5)));
  assign nand_35_nl = ~(main_stage_v_3 & nor_8_cse);
  assign or_179_nl = (fsm_output[0]) | (fsm_output[5]);
  assign nl_AES128_EN_run_staller_inst_run_flen_unreg = MUX1HOT_s_1_5_2(nor_1_nl,
      nor_3_nl, nand_33_nl, nand_34_nl, nand_35_nl, {or_179_nl , (fsm_output[1])
      , (fsm_output[2]) , (fsm_output[3]) , (fsm_output[4])});
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_12_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_12_rg_addr[7:0]),
      .data_out(data_out_out),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_11_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_11_rg_addr[7:0]),
      .data_out(data_out_out_1),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_7_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_7_rg_addr[7:0]),
      .data_out(data_out_out_2),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_1_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_1_rg_addr[7:0]),
      .data_out(data_out_out_3),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_15_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_15_rg_addr[7:0]),
      .data_out(data_out_out_4),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_10_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_10_rg_addr[7:0]),
      .data_out(data_out_out_5),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_rg_addr[7:0]),
      .data_out(data_out_out_6),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_14_rg
      (
      .addr(nl_AES128_EN_SubBytes_1_for_for_read_rom_sbox_rom_map_1_14_rg_addr[7:0]),
      .data_out(data_out_out_7),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_rg
      (
      .addr(nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_rg_addr[7:0]),
      .data_out(data_out_out_8),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_10_rg
      (
      .addr(nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_10_rg_addr[7:0]),
      .data_out(data_out_out_9),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_18_256_8_1  AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_1_rg
      (
      .addr(nl_AES128_EN_SubBytes_for_for_read_rom_sbox_rom_map_1_1_rg_addr[7:0]),
      .data_out(data_out_out_10),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_rg_addr[8:0]),
      .data_out(data_out_out_11),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_14_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_14_rg_addr[8:0]),
      .data_out(data_out_out_12),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_rg_addr[8:0]),
      .data_out(data_out_out_13),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_15_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_15_rg_addr[8:0]),
      .data_out(data_out_out_14),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_11_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_11_rg_addr[8:0]),
      .data_out(data_out_out_15),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_23_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_23_rg_addr[8:0]),
      .data_out(data_out_out_16),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_rg_addr[8:0]),
      .data_out(data_out_out_17),.VDD(VDD),
.VSS(VSS)
    );
  AES128_ENmgc_rom_19_512_8_1  AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_13_rg
      (
      .addr(nl_AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_13_rg_addr[8:0]),
      .data_out(data_out_out_18),.VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_plaintext_in_rsci AES128_EN_run_plaintext_in_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .plaintext_in_rsc_dat(plaintext_in_rsc_dat),
      .plaintext_in_rsc_vld(plaintext_in_rsc_vld),
      .plaintext_in_rsc_rdy(plaintext_in_rsc_rdy),
      .run_wen(run_wen),
      .plaintext_in_rsci_oswt_unreg(or_tmp_49),
      .plaintext_in_rsci_bawt(plaintext_in_rsci_bawt),
      .plaintext_in_rsci_iden(plaintext_in_rsci_iden),
      .plaintext_in_rsci_iswt0(reg_key_in_rsci_iswt0_cse),
      .plaintext_in_rsci_wen_comp(plaintext_in_rsci_wen_comp),
      .plaintext_in_rsci_idat_mxwt(plaintext_in_rsci_idat_mxwt),.VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_key_in_rsci AES128_EN_run_key_in_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .key_in_rsc_dat(key_in_rsc_dat),
      .key_in_rsc_vld(key_in_rsc_vld),
      .key_in_rsc_rdy(key_in_rsc_rdy),
      .run_wen(run_wen),
      .key_in_rsci_oswt_unreg(or_tmp_49),
      .key_in_rsci_bawt(key_in_rsci_bawt),
      .key_in_rsci_iden(key_in_rsci_iden),
      .key_in_rsci_iswt0(reg_key_in_rsci_iswt0_cse),
      .key_in_rsci_wen_comp(key_in_rsci_wen_comp),
      .key_in_rsci_idat_mxwt(key_in_rsci_idat_mxwt),.VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_ciphertext_out_rsci AES128_EN_run_ciphertext_out_rsci_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .ciphertext_out_rsc_dat(ciphertext_out_rsc_dat),
      .ciphertext_out_rsc_vld(ciphertext_out_rsc_vld),
      .ciphertext_out_rsc_rdy(ciphertext_out_rsc_rdy),
      .run_wen(run_wen),
      .ciphertext_out_rsci_oswt_unreg(or_tmp_55),
      .ciphertext_out_rsci_bawt(ciphertext_out_rsci_bawt),
      .ciphertext_out_rsci_iden(ciphertext_out_rsci_iden),
      .ciphertext_out_rsci_iswt0(ciphertext_out_rsci_iswt0),
      .ciphertext_out_rsci_wen_comp(ciphertext_out_rsci_wen_comp),
      .ciphertext_out_rsci_idat(nl_AES128_EN_run_ciphertext_out_rsci_inst_ciphertext_out_rsci_idat[127:0]),.VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_staller AES128_EN_run_staller_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .plaintext_in_rsci_iden(plaintext_in_rsci_iden),
      .plaintext_in_rsci_wen_comp(plaintext_in_rsci_wen_comp),
      .key_in_rsci_iden(key_in_rsci_iden),
      .key_in_rsci_wen_comp(key_in_rsci_wen_comp),
      .ciphertext_out_rsci_iden(ciphertext_out_rsci_iden),
      .ciphertext_out_rsci_wen_comp(ciphertext_out_rsci_wen_comp),
      .run_flen_unreg(nl_AES128_EN_run_staller_inst_run_flen_unreg),.VDD(VDD),
.VSS(VSS)
    );
  AES128_EN_run_run_fsm AES128_EN_run_run_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),.VDD(VDD),
.VSS(VSS)
    );
  assign or_cse = ciphertext_out_rsci_bawt | (~ ROUND_not_mdf_sva_st_1);
  assign and_10_cse = main_stage_v_4 & (~ main_stage_v_5);
  assign nor_8_cse = ~(main_stage_v_4 | main_stage_v_5);
  assign and_546_cse = run_wen & (~((~ (fsm_output[5])) | or_dcpl_67 | (~ ROUND_not_mdf_sva_st)));
  assign ROUND_r_and_cse = run_wen & (~(or_dcpl_66 | or_tmp_118));
  assign or_139_nl = or_tmp_19 | main_stage_v_3 | main_stage_v_1 | (~ main_stage_v_2);
  assign AES128_EN_GenRoundKey_for_mux_33_nl = MUX_s_1_2_2(or_dcpl_49, or_139_nl,
      fsm_output[3]);
  assign AES128_EN_GenRoundKey_for_and_cse = run_wen & (~(AES128_EN_GenRoundKey_for_mux_33_nl
      | or_dcpl_83 | (fsm_output[4])));
  assign state_arr_and_2_cse = run_wen & (~(main_stage_v_4 | (~ main_stage_v_3)))
      & (fsm_output[4]);
  assign state_arr_and_3_cse = run_wen & (~ or_dcpl_90) & (fsm_output[3]);
  assign state_arr_and_4_cse = run_wen & (~ or_dcpl_80) & (fsm_output[3]);
  assign or_145_nl = (~ main_stage_v_4) | main_stage_v_1 | main_stage_v_2;
  assign roundkeys_mux_nl = MUX_s_1_2_2(or_dcpl_49, or_145_nl, fsm_output[5]);
  assign roundkeys_and_cse = run_wen & (~(roundkeys_mux_nl | and_110_cse));
  assign AES128_EN_ShiftRows_a_arr_and_cse = run_wen & (~(or_dcpl | main_stage_v_2))
      & (fsm_output[2]);
  assign AES128_EN_ShiftRows_a_arr_and_1_cse = run_wen & (~(or_dcpl | or_tmp | or_tmp_118));
  assign AES128_EN_MixColumns_for_for_for_else_and_1_cse = run_wen & (~ main_stage_v_2)
      & (fsm_output[2]);
  assign or_134_nl = or_tmp_19 | or_dcpl_80;
  assign AES128_EN_MixColumns_for_for_for_else_mux_18_nl = MUX_s_1_2_2(or_dcpl_76,
      or_134_nl, fsm_output[3]);
  assign AES128_EN_MixColumns_for_for_for_else_and_2_cse = run_wen & (~(AES128_EN_MixColumns_for_for_for_else_mux_18_nl
      | (fsm_output[5]) | (fsm_output[1]) | (fsm_output[4])));
  assign or_164_nl = or_dcpl_110 | or_tmp;
  assign AES128_EN_ShiftRows_a_arr_mux_29_nl = MUX_s_1_2_2(or_dcpl_66, or_164_nl,
      fsm_output[5]);
  assign AES128_EN_ShiftRows_a_arr_and_11_cse = run_wen & (~(AES128_EN_ShiftRows_a_arr_mux_29_nl
      | and_110_cse));
  assign ROUND_and_2_cse = run_wen & (~((~(and_dcpl_36 | and_20_cse)) | or_tmp_118));
  assign AES128_EN_MixColumns_for_for_for_else_and_7_cse = run_wen & (~(main_stage_v_1
      | or_tmp_118));
  assign ROUND_and_9_cse = run_wen & (~((~(and_dcpl_35 | and_dcpl)) | or_tmp_118));
  assign AES128_EN_AddRoundKey_2_for_for_and_cse = run_wen & (~ or_dcpl) & (fsm_output[3]);
  assign AES128_EN_GenRoundKey_1_for_and_cse = run_wen & (~ main_stage_v_3) & (fsm_output[3]);
  assign and_20_cse = and_dcpl & (~ main_stage_v_2);
  assign AES128_EN_AddRoundKey_2_for_for_and_15_cse = run_wen & (~ main_stage_v_4)
      & (fsm_output[4]);
  assign ROUND_ROUND_and_tmp = (ROUND_r_3_0_sva_2[3:1]==3'b101);
  assign nl_ROUND_r_3_0_sva_2 = ROUND_r_3_0_lpi_1_dfm_mx0 + 4'b0001;
  assign ROUND_r_3_0_sva_2 = nl_ROUND_r_3_0_sva_2[3:0];
  assign AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1 =
      AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva ^ data_out_out_8
      ^ AES128_EN_Rcon_mux_itm;
  assign state_arr_3_1_1_sva_2 = data_out_out_16 ^ AES128_EN_ShiftRows_a_arr_1_1_sva
      ^ AES128_EN_ShiftRows_a_arr_2_1_sva ^ data_out_out_14 ^ AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  assign state_arr_3_0_1_sva_2 = AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_8_itm
      ^ AES128_EN_ShiftRows_a_arr_1_0_sva ^ AES128_EN_ShiftRows_a_arr_2_0_sva ^ data_out_out_13
      ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
  assign state_arr_1_1_1_sva_2 = AES128_EN_ShiftRows_a_arr_0_1_sva ^ data_out_out_13
      ^ data_out_out_16 ^ AES128_EN_ShiftRows_a_arr_3_1_sva ^ AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  assign state_arr_1_2_1_sva_2 = AES128_EN_ShiftRows_a_arr_0_2_sva ^ data_out_out_18
      ^ data_out_out_11 ^ AES128_EN_ShiftRows_a_arr_3_2_sva ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  assign state_arr_2_3_1_sva_2 = AES128_EN_ShiftRows_a_arr_0_3_sva ^ AES128_EN_ShiftRows_a_arr_1_3_sva
      ^ data_out_out_17 ^ data_out_out_15 ^ AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  assign state_arr_2_2_1_sva_2 = AES128_EN_ShiftRows_a_arr_0_2_sva ^ AES128_EN_ShiftRows_a_arr_1_2_sva
      ^ data_out_out_11 ^ data_out_out_18 ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
  assign main_stage_v_5_mx1 = main_stage_v_5 & ROUND_not_mdf_sva_st_1 & (~ ciphertext_out_rsci_bawt);
  assign ROUND_r_3_0_lpi_1_dfm_mx0 = MUX_v_4_2_2(ROUND_r_3_0_sva_1, 4'b0001, exitL_exit_ROUND_sva);
  assign or_dcpl = main_stage_v_4 | main_stage_v_3;
  assign and_dcpl = ~(exitL_exit_ROUND_sva | main_stage_v_1);
  assign or_tmp = main_stage_v_2 | main_stage_v_1;
  assign nor_17_cse = ~(main_stage_v_1 | main_stage_v_2);
  assign or_tmp_19 = main_stage_v_4 | main_stage_v_5;
  assign and_dcpl_35 = exitL_exit_ROUND_sva & (~ main_stage_v_1);
  assign and_dcpl_36 = and_dcpl_35 & (~ main_stage_v_2);
  assign or_dcpl_43 = ~(main_stage_v_5 & main_stage_v_4);
  assign or_dcpl_45 = (~(main_stage_v_5 & ROUND_not_mdf_sva_st_1)) | ciphertext_out_rsci_bawt;
  assign or_dcpl_48 = (~ exitL_exit_ROUND_sva) | main_stage_v_1;
  assign or_dcpl_49 = or_dcpl_48 | main_stage_v_2;
  assign and_dcpl_49 = main_stage_v_5 & ROUND_not_mdf_sva_st_1;
  assign nand_26_cse = ~(key_in_rsci_bawt & plaintext_in_rsci_bawt);
  assign or_dcpl_66 = (and_dcpl_49 & (~ ciphertext_out_rsci_bawt)) | (nand_26_cse
      & ROUND_asn_itm) | (~ main_stage_v) | main_stage_v_4 | main_stage_v_3 | or_tmp;
  assign or_dcpl_67 = main_stage_v_5 | (~ main_stage_v_4);
  assign or_dcpl_76 = (~ main_stage_v_1) | main_stage_v_2;
  assign or_dcpl_80 = main_stage_v_3 | (~ main_stage_v_2);
  assign or_dcpl_83 = (fsm_output[5]) | (fsm_output[2]);
  assign or_dcpl_88 = or_dcpl | or_dcpl_76;
  assign or_dcpl_90 = or_dcpl | (~ main_stage_v_2);
  assign or_dcpl_94 = (~ main_stage_v_3) | main_stage_v_1;
  assign or_dcpl_110 = or_dcpl_67 | main_stage_v_3;
  assign or_tmp_49 = or_dcpl_45 & main_stage_v & key_in_rsci_bawt & plaintext_in_rsci_bawt
      & ROUND_asn_itm & (~ main_stage_v_4) & (~ main_stage_v_3) & nor_17_cse & (fsm_output[1]);
  assign and_110_cse = (fsm_output[4:2]!=3'b000);
  assign or_tmp_55 = and_dcpl_49 & ciphertext_out_rsci_bawt & (fsm_output[1]);
  assign or_tmp_98 = (~(nand_26_cse & ROUND_asn_itm)) & or_dcpl_45 & main_stage_v
      & (~ main_stage_v_4) & (~ main_stage_v_3) & nor_17_cse & (fsm_output[1]);
  assign or_tmp_99 = or_dcpl_43 & (~ main_stage_v) & (~(main_stage_v_3 | main_stage_v_1
      | main_stage_v_2)) & (fsm_output[5]);
  assign or_tmp_103 = nor_8_cse & (~ main_stage_v_3) & main_stage_v_1 & (~ main_stage_v_2)
      & (fsm_output[2]);
  assign or_tmp_107 = nor_8_cse & (~ main_stage_v_3) & main_stage_v_2 & (fsm_output[3]);
  assign or_tmp_111 = nor_8_cse & main_stage_v_3 & (fsm_output[4]);
  assign or_tmp_115 = and_10_cse & (fsm_output[5]);
  assign or_tmp_118 = ~((fsm_output[1:0]!=2'b00));
  assign or_tmp_145 = or_dcpl_83 | (fsm_output[3]);
  assign main_stage_v_5_mx0c0 = or_cse & main_stage_v_5 & (fsm_output[1]);
  assign xor_cse = AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva
      ^ data_out_out_8 ^ AES128_EN_Rcon_mux_itm ^ AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  assign AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1 =
      AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva ^ xor_cse;
  assign state_arr_0_1_1_sva_2 = xor_cse ^ data_out_out_17 ^ data_out_out_13 ^ AES128_EN_ShiftRows_a_arr_2_1_sva
      ^ AES128_EN_ShiftRows_a_arr_3_1_sva;
  assign state_arr_0_2_1_sva_2 = AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva
      ^ xor_cse ^ data_out_out_16 ^ data_out_out_18 ^ AES128_EN_ShiftRows_a_arr_2_2_sva
      ^ AES128_EN_ShiftRows_a_arr_3_2_sva;
  assign state_arr_0_3_1_sva_2 = xor_cse ^ data_out_out_14 ^ data_out_out_15 ^ AES128_EN_ShiftRows_a_arr_2_3_sva
      ^ AES128_EN_ShiftRows_a_arr_3_3_sva ^ roundkeys_12_lpi_1 ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva;
  assign xor_cse_14 = MUX_v_8_2_2(AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_7_ncse_sva,
      (key_in_rsci_idat_mxwt[39:32]), exitL_exit_ROUND_sva);
  assign xor_cse_15 = MUX_v_8_2_2(AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva,
      (key_in_rsci_idat_mxwt[71:64]), exitL_exit_ROUND_sva);
  assign xor_cse_16 = MUX_v_8_2_2(AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva,
      (key_in_rsci_idat_mxwt[103:96]), exitL_exit_ROUND_sva);
  assign for_1_mux_8_nl = MUX_v_8_2_2(roundkeys_15_lpi_1, (key_in_rsci_idat_mxwt[7:0]),
      exitL_exit_ROUND_sva);
  assign xor_cse_13 = xor_cse_14 ^ xor_cse_15 ^ xor_cse_16 ^ for_1_mux_8_nl;
  assign xor_cse_22 = ROUND_mux_10_itm ^ ROUND_mux_6_itm ^ ROUND_mux_2_itm ^ roundkeys_13_lpi_1;
  assign xor_cse_27 = (AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[0])
      ^ (xor_cse[0]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[0]);
  assign xor_cse_34 = (AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[2:1])
      ^ (xor_cse[2:1]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[2:1]);
  assign xor_cse_41 = (AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[3])
      ^ (xor_cse[3]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[3]);
  assign xor_cse_48 = (AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[5:4])
      ^ (xor_cse[5:4]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[5:4]);
  assign xor_cse_55 = (AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[7:6])
      ^ (xor_cse[7:6]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[7:6]);
  assign AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0
      = roundkeys_12_lpi_1 ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva
      ^ xor_cse;
  assign AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva_mx1w0
      = data_out_out_9 ^ xor_cse_22;
  assign xor_cse_69 = ROUND_mux_3_itm ^ data_out_out_2 ^ ROUND_mux_11_itm;
  assign xor_cse_72 = AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva
      ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_3_ncse_sva ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
  assign AES128_EN_MixColumns_for_for_for_else_nor_1_cse = ~((fsm_output[5]) | (fsm_output[3]));
  assign AES128_EN_SubBytes_1_for_for_and_cse = (~ exitL_exit_ROUND_sva) & (fsm_output[1]);
  assign AES128_EN_SubBytes_1_for_for_and_1_cse = exitL_exit_ROUND_sva & (fsm_output[1]);
  assign AES128_EN_MixColumns_for_for_for_else_or_cse = (fsm_output[2:1]!=2'b00);
  assign AES128_EN_MixColumns_for_for_for_else_or_1_cse = (fsm_output[5:4]!=2'b00);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_key_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( rst ) begin
      reg_key_in_rsci_iswt0_cse <= 1'b0;
    end
    else if ( run_wen & ((or_dcpl_43 & (~(main_stage_v | main_stage_v_3)) & and_dcpl_36
        & (fsm_output[5])) | (fsm_output[0]) | or_tmp_49) ) begin
      reg_key_in_rsci_iswt0_cse <= ~ or_tmp_49;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      exitL_exit_ROUND_sva <= 1'b1;
    end
    else if ( rst ) begin
      exitL_exit_ROUND_sva <= 1'b1;
    end
    else if ( run_wen & (~((~ (fsm_output[1])) | or_dcpl_66)) ) begin
      exitL_exit_ROUND_sva <= ROUND_ROUND_and_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ciphertext_out_rsci_iswt0 <= 1'b0;
    end
    else if ( rst ) begin
      ciphertext_out_rsci_iswt0 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_55 | (and_10_cse & ROUND_not_mdf_sva_st & (fsm_output[5])))
        ) begin
      ciphertext_out_rsci_iswt0 <= ~ or_tmp_55;
    end
  end
  always @(posedge clk) begin
    if ( and_546_cse ) begin
      ciphertext_out_rsci_idat_59 <= AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_61_60 <= AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
      ciphertext_out_rsci_idat_58_57 <= AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
      ciphertext_out_rsci_idat_63_62 <= AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
      ciphertext_out_rsci_idat_56 <= AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
      ciphertext_out_rsci_idat_71_64 <= data_out_out ^ AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva;
      ciphertext_out_rsci_idat_55_48 <= AES128_EN_AddRoundKey_2_for_2_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_79_72 <= data_out_out_1 ^ AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
      ciphertext_out_rsci_idat_47_40 <= data_out_out_2 ^ AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
      ciphertext_out_rsci_idat_87_80 <= AES128_EN_AddRoundKey_2_for_2_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_39_32 <= data_out_out_3 ^ AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva;
      ciphertext_out_rsci_idat_88 <= AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
      ciphertext_out_rsci_idat_31_30 <= AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
      ciphertext_out_rsci_idat_90_89 <= AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
      ciphertext_out_rsci_idat_29_28 <= AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
      ciphertext_out_rsci_idat_91 <= AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_27 <= AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_93_92 <= AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_3_itm;
      ciphertext_out_rsci_idat_26_25 <= AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_2_itm;
      ciphertext_out_rsci_idat_95_94 <= AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_5_itm;
      ciphertext_out_rsci_idat_24 <= AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_4_itm;
      ciphertext_out_rsci_idat_103_96 <= AES128_EN_AddRoundKey_2_for_4_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_23_16 <= data_out_out_4 ^ AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva
          ^ AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_3_ncse_sva;
      ciphertext_out_rsci_idat_111_104 <= data_out_out_5 ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
      ciphertext_out_rsci_idat_15_8 <= data_out_out_6 ^ AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva
          ^ AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva;
      ciphertext_out_rsci_idat_119_112 <= AES128_EN_AddRoundKey_2_for_2_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm;
      ciphertext_out_rsci_idat_7_0 <= data_out_out_7 ^ AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_7_ncse_sva
          ^ AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva;
      ciphertext_out_rsci_idat_123 <= AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_3;
      ciphertext_out_rsci_idat_122_121 <= AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_2_1;
      ciphertext_out_rsci_idat_125_124 <= AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_5_4;
      ciphertext_out_rsci_idat_120 <= AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_0;
      ciphertext_out_rsci_idat_127_126 <= AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_7_6;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v <= 1'b1;
    end
    else if ( rst ) begin
      main_stage_v <= 1'b1;
    end
    else if ( run_wen & (or_tmp_98 | or_tmp_99) ) begin
      main_stage_v <= ~ or_tmp_98;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_98 | or_tmp_103) ) begin
      main_stage_v_1 <= ~ or_tmp_103;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_103 | or_tmp_107) ) begin
      main_stage_v_2 <= ~ or_tmp_107;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_107 | or_tmp_111) ) begin
      main_stage_v_3 <= ~ or_tmp_111;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( run_wen & (or_tmp_111 | or_tmp_115) ) begin
      main_stage_v_4 <= ~ or_tmp_115;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROUND_asn_itm <= 1'b1;
    end
    else if ( rst ) begin
      ROUND_asn_itm <= 1'b1;
    end
    else if ( run_wen & or_tmp_99 ) begin
      ROUND_asn_itm <= exitL_exit_ROUND_sva;
    end
  end
  always @(posedge clk) begin
    if ( ROUND_r_and_cse ) begin
      ROUND_r_3_0_sva_1 <= ROUND_r_3_0_sva_2;
      state_arr_3_3_1_lpi_1 <= data_out_out_6 ^ xor_cse_13 ^ data_out_out_11 ^ data_out_out_5
          ^ data_out_out_4 ^ data_out_out_12;
      AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_7_ncse_sva <= xor_cse_14
          ^ xor_cse_15 ^ xor_cse_16 ^ data_out_out_6;
      AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva <= xor_cse_15
          ^ xor_cse_16 ^ data_out_out_6;
      AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva <= xor_cse_16
          ^ data_out_out_6;
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_GenRoundKey_for_and_cse ) begin
      AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[63:56]),
          AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1,
          fsm_output[3]);
      AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_1_ncse_sva <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[95:88]),
          xor_cse, fsm_output[3]);
      AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[127:120]),
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1,
          fsm_output[3]);
      ROUND_mux_20_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_1_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          state_arr_0_1_1_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~ or_dcpl_88) & (fsm_output[2]) ) begin
      state_arr_3_2_1_lpi_1 <= AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_4_itm
          ^ data_out_out_7 ^ AES128_EN_ShiftRows_a_arr_2_2_sva ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_5_itm
          ^ AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_7_ncse_sva;
    end
  end
  always @(posedge clk) begin
    if ( state_arr_and_2_cse ) begin
      state_arr_2_1_1_lpi_1 <= AES128_EN_ShiftRows_a_arr_0_1_sva ^ AES128_EN_ShiftRows_a_arr_1_1_sva
          ^ data_out_out_12 ^ data_out_out_14 ^ AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva;
      state_arr_1_0_1_lpi_1 <= AES128_EN_ShiftRows_a_arr_0_0_sva ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_24_itm
          ^ data_out_out_15 ^ AES128_EN_ShiftRows_a_arr_3_0_sva ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva;
    end
  end
  always @(posedge clk) begin
    if ( state_arr_and_3_cse ) begin
      state_arr_2_0_1_lpi_1 <= AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_16_itm
          ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_itm
          ^ AES128_EN_ShiftRows_a_arr_0_0_sva ^ AES128_EN_ShiftRows_a_arr_1_0_sva
          ^ ROUND_mux_3_itm ^ data_out_out_2;
      AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_5_ncse_sva <= ROUND_mux_7_itm
          ^ xor_cse_69;
    end
  end
  always @(posedge clk) begin
    if ( state_arr_and_4_cse ) begin
      state_arr_1_3_1_lpi_1 <= data_out_out_9 ^ xor_cse_22 ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_18_itm
          ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_19_itm
          ^ AES128_EN_ShiftRows_a_arr_0_3_sva ^ AES128_EN_ShiftRows_a_arr_3_3_sva;
      state_arr_0_0_lpi_1 <= AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_itm
          ^ AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_itm
          ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva
          ^ data_out_out_8 ^ AES128_EN_Rcon_mux_itm ^ AES128_EN_ShiftRows_a_arr_2_0_sva
          ^ AES128_EN_ShiftRows_a_arr_3_0_sva;
      AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva <= ROUND_mux_3_itm
          ^ data_out_out_2;
      AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_3_ncse_sva <= ROUND_mux_10_itm
          ^ ROUND_mux_6_itm ^ ROUND_mux_2_itm ^ data_out_out_9;
      AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva <= ROUND_mux_7_itm
          ^ ROUND_mux_3_itm ^ data_out_out_2;
      AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva <= ROUND_mux_6_itm
          ^ ROUND_mux_2_itm ^ data_out_out_9;
      AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva <= ROUND_mux_2_itm
          ^ data_out_out_9;
    end
  end
  always @(posedge clk) begin
    if ( roundkeys_and_cse ) begin
      roundkeys_15_lpi_1 <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[7:0]), AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_7_ncse_sva,
          fsm_output[5]);
      roundkeys_14_lpi_1 <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[15:8]), AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva,
          fsm_output[5]);
      roundkeys_13_lpi_1 <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[23:16]), AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva,
          fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(roundkeys_mux_3_nl | or_tmp_145)) ) begin
      roundkeys_12_lpi_1 <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[31:24]), AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva,
          fsm_output[4]);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_ShiftRows_a_arr_and_cse ) begin
      AES128_EN_ShiftRows_a_arr_1_2_sva <= data_out_out_7;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_8_itm
          <= data_out_out_16;
      AES128_EN_ShiftRows_a_arr_3_0_sva <= data_out_out_2;
      AES128_EN_ShiftRows_a_arr_2_0_sva <= data_out_out_9;
      AES128_EN_ShiftRows_a_arr_3_1_sva <= data_out_out_4;
      AES128_EN_ShiftRows_a_arr_1_1_sva <= data_out_out_6;
      AES128_EN_ShiftRows_a_arr_2_1_sva <= data_out_out_5;
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_ShiftRows_a_arr_and_1_cse ) begin
      AES128_EN_ShiftRows_a_arr_2_2_sva <= data_out_out_7;
      AES128_EN_ShiftRows_a_arr_2_3_sva <= data_out_out_4;
      AES128_EN_ShiftRows_a_arr_1_3_sva <= data_out_out_5;
      AES128_EN_ShiftRows_a_arr_3_3_sva <= data_out_out_9;
      AES128_EN_ShiftRows_a_arr_3_2_sva <= data_out_out_2;
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_7_ncse_sva <= data_out_out_6
          ^ xor_cse_13;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(AES128_EN_ShiftRows_a_arr_mux_27_nl | (fsm_output[5]) | (fsm_output[3])
        | (fsm_output[1]))) ) begin
      AES128_EN_ShiftRows_a_arr_0_0_sva <= MUX_v_8_2_2(data_out_out_8, state_arr_1_1_1_sva_2,
          fsm_output[4]);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_MixColumns_for_for_for_else_and_1_cse ) begin
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_17_itm
          <= data_out_out_13;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_19_itm
          <= data_out_out_14;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_18_itm
          <= data_out_out_15;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_itm <=
          data_out_out_11;
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_MixColumns_for_for_for_else_and_2_cse ) begin
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_16_itm
          <= MUX_v_8_2_2(data_out_out_12, state_arr_0_3_1_sva_2, fsm_output[3]);
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_1_itm
          <= MUX_v_8_2_2(data_out_out_17, state_arr_0_2_1_sva_2, fsm_output[3]);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(AES128_EN_ShiftRows_a_arr_mux_28_nl | (fsm_output[3]) | (fsm_output[1])
        | (fsm_output[4]))) ) begin
      AES128_EN_ShiftRows_a_arr_1_0_sva <= MUX_v_8_2_2(data_out_out_10, state_arr_3_1_1_sva_2,
          fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_ShiftRows_a_arr_and_11_cse ) begin
      AES128_EN_ShiftRows_a_arr_0_3_sva <= MUX_v_8_2_2(data_out_out_10, state_arr_3_0_1_sva_2,
          fsm_output[5]);
      AES128_EN_ShiftRows_a_arr_0_2_sva <= MUX_v_8_2_2(data_out_out_8, state_arr_2_3_1_sva_2,
          fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( ROUND_and_2_cse ) begin
      ROUND_mux_11_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[47:40]), AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_5_ncse_sva,
          and_20_cse);
      ROUND_mux_10_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[55:48]), AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_3_ncse_sva,
          and_20_cse);
      ROUND_mux_7_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[79:72]), AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva,
          and_20_cse);
      ROUND_mux_6_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[87:80]), AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva,
          and_20_cse);
      ROUND_mux_3_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[111:104]), AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva,
          and_20_cse);
      ROUND_mux_2_itm <= MUX_v_8_2_2((key_in_rsci_idat_mxwt[119:112]), AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva,
          and_20_cse);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(or_tmp | or_tmp_118)) ) begin
      AES128_EN_Rcon_mux_itm <= MUX_v_8_10_2x0(8'b00000001, 8'b00000010, 8'b00000100,
          8'b00001000, 8'b00010000, 8'b00100000, 8'b01000000, 8'b10000000, 8'b00011011,
          ROUND_r_3_0_lpi_1_dfm_mx0);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_MixColumns_for_for_for_else_and_7_cse ) begin
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_4_itm
          <= data_out_out_16;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_5_itm
          <= data_out_out_13;
    end
  end
  always @(posedge clk) begin
    if ( ROUND_and_9_cse ) begin
      ROUND_mux_31_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_4_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          AES128_EN_ShiftRows_a_arr_0_3_sva, and_dcpl);
      ROUND_mux_34_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_4_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          state_arr_3_3_1_lpi_1, and_dcpl);
      ROUND_mux_24_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_2_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          AES128_EN_ShiftRows_a_arr_0_0_sva, and_dcpl);
      ROUND_mux_26_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_2_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          state_arr_1_3_1_lpi_1, and_dcpl);
      ROUND_mux_30_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_3_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          AES128_EN_ShiftRows_a_arr_0_2_sva, and_dcpl);
      ROUND_mux_29_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_3_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          AES128_EN_ShiftRows_a_arr_0_1_sva, and_dcpl);
      ROUND_mux_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_1_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          state_arr_0_0_lpi_1, and_dcpl);
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(ROUND_mux_53_nl | or_tmp_145)) ) begin
      ROUND_mux_25_itm <= MUX_v_8_2_2(AES128_EN_AddRoundKey_for_2_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl,
          state_arr_1_2_1_sva_2, fsm_output[4]);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_AddRoundKey_2_for_for_and_cse ) begin
      AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_4_itm
          <= (data_out_out_1[0]) ^ (AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0[0])
          ^ (data_out_out_5[0]) ^ xor_cse_27;
      AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_2_itm
          <= ~((data_out_out_1[2:1]) ^ (AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0[2:1])
          ^ (data_out_out_5[2:1]) ^ xor_cse_34);
      AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= (data_out_out_1[3]) ^ (AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0[3])
          ^ (data_out_out_5[3]) ^ xor_cse_41;
      AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_3_itm
          <= ~((data_out_out_1[5:4]) ^ (AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0[5:4])
          ^ (data_out_out_5[5:4]) ^ xor_cse_48);
      AES128_EN_AddRoundKey_2_for_1_for_4_AES128_EN_AddRoundKey_2_for_for_xor_5_itm
          <= (data_out_out_1[7:6]) ^ (AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0[7:6])
          ^ (data_out_out_5[7:6]) ^ xor_cse_55;
      AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_4_itm
          <= (data_out_out[0]) ^ (data_out_out_5[0]) ^ xor_cse_27;
      AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_2_itm
          <= ~((data_out_out[2:1]) ^ (data_out_out_5[2:1]) ^ xor_cse_34);
      AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= (data_out_out[3]) ^ (data_out_out_5[3]) ^ xor_cse_41;
      AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_3_itm
          <= ~((data_out_out[5:4]) ^ (data_out_out_5[5:4]) ^ xor_cse_48);
      AES128_EN_AddRoundKey_2_for_1_for_3_AES128_EN_AddRoundKey_2_for_for_xor_5_itm
          <= (data_out_out[7:6]) ^ (data_out_out_5[7:6]) ^ xor_cse_55;
      AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_4_itm
          <= (data_out_out_3[0]) ^ (xor_cse[0]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[0])
          ^ (data_out_out_5[0]);
      AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_2_itm
          <= ~((data_out_out_3[2:1]) ^ (xor_cse[2:1]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[2:1])
          ^ (data_out_out_5[2:1]));
      AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= (data_out_out_3[3]) ^ (xor_cse[3]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[3])
          ^ (data_out_out_5[3]);
      AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_3_itm
          <= ~((data_out_out_3[5:4]) ^ (xor_cse[5:4]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[5:4])
          ^ (data_out_out_5[5:4]));
      AES128_EN_AddRoundKey_2_for_1_for_2_AES128_EN_AddRoundKey_2_for_for_xor_5_itm
          <= (data_out_out_3[7:6]) ^ (xor_cse[7:6]) ^ (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[7:6])
          ^ (data_out_out_5[7:6]);
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva <= AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_3_ncse_sva_mx1w0;
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_5_ncse_sva <= roundkeys_14_lpi_1
          ^ ROUND_mux_7_itm ^ xor_cse_69;
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_GenRoundKey_1_for_and_cse ) begin
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_7_6_sva
          <= (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[7:6])
          ^ (data_out_out_5[7:6]);
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_0_sva
          <= (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[0])
          ^ (data_out_out_5[0]);
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_5_4_sva
          <= ~((AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[5:4])
          ^ (data_out_out_5[5:4]));
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_2_1_sva
          <= ~((AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[2:1])
          ^ (data_out_out_5[2:1]));
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_3_sva
          <= (AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_1[3])
          ^ (data_out_out_5[3]);
      AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva <= AES128_EN_GenRoundKey_for_4_AES128_EN_GenRoundKey_for_xor_1_ncse_sva_mx1w0;
      AES128_EN_MixColumns_for_for_for_else_read_rom_GF_MUL_TABLE_rom_map_1_24_itm
          <= data_out_out_12;
    end
  end
  always @(posedge clk) begin
    if ( run_wen & (~(AES128_EN_ShiftRows_a_arr_mux_31_nl | (fsm_output[2]) | (fsm_output[1])
        | (fsm_output[4]))) ) begin
      AES128_EN_ShiftRows_a_arr_0_1_sva <= MUX_v_8_2_2(data_out_out_10, state_arr_2_2_1_sva_2,
          fsm_output[5]);
    end
  end
  always @(posedge clk) begin
    if ( AES128_EN_AddRoundKey_2_for_for_and_15_cse ) begin
      AES128_EN_AddRoundKey_2_for_2_for_3_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= data_out_out_2 ^ data_out_out_9 ^ xor_cse_72;
      AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_3_ncse_sva <=
          data_out_out_9 ^ xor_cse_72;
      AES128_EN_AddRoundKey_2_for_2_for_2_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= data_out_out ^ AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_3_ncse_sva
          ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva
          ^ data_out_out_9;
      AES128_EN_AddRoundKey_2_for_4_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= data_out_out_4 ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva
          ^ data_out_out_5;
      AES128_EN_AddRoundKey_2_for_2_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm
          <= data_out_out_3 ^ AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_3_ncse_sva
          ^ data_out_out_9;
      AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_7_6
          <= (data_out_out_6[7:6]) ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_7_6_sva;
      AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_0
          <= (data_out_out_6[0]) ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_0_sva;
      AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_5_4
          <= (data_out_out_6[5:4]) ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_5_4_sva;
      AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_2_1
          <= (data_out_out_6[2:1]) ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_2_1_sva;
      AES128_EN_AddRoundKey_2_for_1_for_1_AES128_EN_AddRoundKey_2_for_for_xor_1_itm_3
          <= (data_out_out_6[3]) ^ AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_1_ncse_3_sva;
      AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva <=
          AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_7_ncse_sva ^
          AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva ^
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva ^
          data_out_out_5;
      AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_7_ncse_sva <=
          AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_7_ncse_sva ^
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_7_ncse_sva ^
          data_out_out_5;
      AES128_EN_GenRoundKey_1_for_3_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva <=
          AES128_EN_GenRoundKey_for_3_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          data_out_out_7;
      AES128_EN_GenRoundKey_1_for_2_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva <=
          AES128_EN_GenRoundKey_for_2_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          data_out_out_7;
      AES128_EN_GenRoundKey_1_for_1_AES128_EN_GenRoundKey_1_for_xor_5_ncse_sva <=
          AES128_EN_GenRoundKey_for_1_AES128_EN_GenRoundKey_for_xor_5_ncse_sva ^
          data_out_out_7;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROUND_not_mdf_sva_st <= 1'b0;
    end
    else if ( rst ) begin
      ROUND_not_mdf_sva_st <= 1'b0;
    end
    else if ( AES128_EN_ShiftRows_a_arr_and_1_cse ) begin
      ROUND_not_mdf_sva_st <= ROUND_ROUND_and_tmp;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( rst ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( run_wen & (main_stage_v_5_mx0c0 | or_tmp_115) ) begin
      main_stage_v_5 <= ~ main_stage_v_5_mx0c0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ROUND_not_mdf_sva_st_1 <= 1'b0;
    end
    else if ( rst ) begin
      ROUND_not_mdf_sva_st_1 <= 1'b0;
    end
    else if ( run_wen & or_tmp_115 ) begin
      ROUND_not_mdf_sva_st_1 <= ROUND_not_mdf_sva_st;
    end
  end
  assign AES128_EN_AddRoundKey_for_1_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[95:88]) ^ (key_in_rsci_idat_mxwt[95:88]);
  assign or_148_nl = or_dcpl_94 | main_stage_v_2;
  assign roundkeys_mux_3_nl = MUX_s_1_2_2(or_dcpl_49, or_148_nl, fsm_output[4]);
  assign or_154_nl = main_stage_v_3 | (~ main_stage_v_1) | main_stage_v_2;
  assign or_156_nl = or_tmp_19 | (~ main_stage_v_3) | main_stage_v_2;
  assign AES128_EN_ShiftRows_a_arr_mux_27_nl = MUX_s_1_2_2(or_154_nl, or_156_nl,
      fsm_output[4]);
  assign or_162_nl = or_dcpl_67 | main_stage_v_3 | main_stage_v_2;
  assign AES128_EN_ShiftRows_a_arr_mux_28_nl = MUX_s_1_2_2(or_dcpl_88, or_162_nl,
      fsm_output[5]);
  assign AES128_EN_AddRoundKey_for_4_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[103:96]) ^ (key_in_rsci_idat_mxwt[103:96]);
  assign AES128_EN_AddRoundKey_for_4_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[7:0]) ^ (key_in_rsci_idat_mxwt[7:0]);
  assign AES128_EN_AddRoundKey_for_2_for_2_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[87:80]) ^ (key_in_rsci_idat_mxwt[87:80]);
  assign AES128_EN_AddRoundKey_for_2_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[23:16]) ^ (key_in_rsci_idat_mxwt[23:16]);
  assign AES128_EN_AddRoundKey_for_3_for_4_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[15:8]) ^ (key_in_rsci_idat_mxwt[15:8]);
  assign AES128_EN_AddRoundKey_for_3_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[47:40]) ^ (key_in_rsci_idat_mxwt[47:40]);
  assign AES128_EN_AddRoundKey_for_1_for_1_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[127:120]) ^ (key_in_rsci_idat_mxwt[127:120]);
  assign AES128_EN_AddRoundKey_for_2_for_3_AES128_EN_AddRoundKey_for_for_xor_1_nl
      = (plaintext_in_rsci_idat_mxwt[55:48]) ^ (key_in_rsci_idat_mxwt[55:48]);
  assign ROUND_mux_53_nl = MUX_s_1_2_2(or_dcpl_48, or_dcpl_94, fsm_output[4]);
  assign AES128_EN_ShiftRows_a_arr_mux_31_nl = MUX_s_1_2_2(or_dcpl_90, or_dcpl_110,
      fsm_output[5]);

  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_3_2;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [2:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    MUX1HOT_v_8_3_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_4_2;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [3:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    MUX1HOT_v_8_4_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_5_2;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [4:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    MUX1HOT_v_8_5_2 = result;
  end
  endfunction


  function automatic [7:0] MUX1HOT_v_8_6_2;
    input [7:0] input_5;
    input [7:0] input_4;
    input [7:0] input_3;
    input [7:0] input_2;
    input [7:0] input_1;
    input [7:0] input_0;
    input [5:0] sel;
    reg [7:0] result;
  begin
    result = input_0 & {8{sel[0]}};
    result = result | (input_1 & {8{sel[1]}});
    result = result | (input_2 & {8{sel[2]}});
    result = result | (input_3 & {8{sel[3]}});
    result = result | (input_4 & {8{sel[4]}});
    result = result | (input_5 & {8{sel[5]}});
    MUX1HOT_v_8_6_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_10_2x0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [7:0] input_8;
    input [7:0] input_9;
    input [3:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      4'b0001 : begin
        result = input_1;
      end
      4'b0010 : begin
        result = input_2;
      end
      4'b0011 : begin
        result = input_3;
      end
      4'b0100 : begin
        result = input_4;
      end
      4'b0101 : begin
        result = input_5;
      end
      4'b0110 : begin
        result = input_6;
      end
      4'b0111 : begin
        result = input_7;
      end
      4'b1000 : begin
        result = input_8;
      end
      default : begin
        result = input_9;
      end
    endcase
    MUX_v_8_10_2x0 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    AES128_EN
// ------------------------------------------------------------------


module AES128_EN (
  clk, rst, arst_n, plaintext_in_rsc_dat, plaintext_in_rsc_vld, plaintext_in_rsc_rdy,
      key_in_rsc_dat, key_in_rsc_vld, key_in_rsc_rdy, ciphertext_out_rsc_dat, ciphertext_out_rsc_vld,
      ciphertext_out_rsc_rdy,.VDD(VDD),
.VSS(VSS)
);
  input clk;
  input rst;
  input arst_n;
  input [127:0] plaintext_in_rsc_dat;
  input plaintext_in_rsc_vld;
  output plaintext_in_rsc_rdy;
  input [127:0] key_in_rsc_dat;
  input key_in_rsc_vld;
  output key_in_rsc_rdy;
  output [127:0] ciphertext_out_rsc_dat;
  output ciphertext_out_rsc_vld;
  input ciphertext_out_rsc_rdy;
  input VDD;
  input VSS;


  // Interconnect Declarations for Component Instantiations 
  AES128_EN_run AES128_EN_run_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .plaintext_in_rsc_dat(plaintext_in_rsc_dat),
      .plaintext_in_rsc_vld(plaintext_in_rsc_vld),
      .plaintext_in_rsc_rdy(plaintext_in_rsc_rdy),
      .key_in_rsc_dat(key_in_rsc_dat),
      .key_in_rsc_vld(key_in_rsc_vld),
      .key_in_rsc_rdy(key_in_rsc_rdy),
      .ciphertext_out_rsc_dat(ciphertext_out_rsc_dat),
      .ciphertext_out_rsc_vld(ciphertext_out_rsc_vld),
      .ciphertext_out_rsc_rdy(ciphertext_out_rsc_rdy),.VDD(VDD),
.VSS(VSS)
    );
endmodule



