
//------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.2/1059873 Production Release
//  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
// 
//  Generated by:   r12016@cad40
//  Generated date: Thu Jun 13 02:36:44 2024
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
// ------------------------------------------------------------------


module UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
    (
  clken, we, d, wadr, clken_d, d_d, wadr_d, we_d, writeA_w_ram_ir_internal_WMASK_B_d
);
  output clken;
  output we;
  output [11:0] d;
  output [14:0] wadr;
  input clken_d;
  input [11:0] d_d;
  input [14:0] wadr_d;
  input we_d;
  input writeA_w_ram_ir_internal_WMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign we = (writeA_w_ram_ir_internal_WMASK_B_d);
  assign d = (d_d);
  assign wadr = (wadr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
// ------------------------------------------------------------------


module UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
    (
  clken, q, re, radr, clken_d, q_d, radr_d, re_d, readA_r_ram_ir_internal_RMASK_B_d
);
  output clken;
  input [11:0] q;
  output re;
  output [14:0] radr;
  input clken_d;
  output [11:0] q_d;
  input [14:0] radr_d;
  input re_d;
  input readA_r_ram_ir_internal_RMASK_B_d;



  // Interconnect Declarations for Component Instantiations 
  assign clken = (clken_d);
  assign q_d = q;
  assign re = (readA_r_ram_ir_internal_RMASK_B_d);
  assign radr = (radr_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    UNET_IP_maxpool_run_max_run_max_fsm
//  FSM Module
// ------------------------------------------------------------------


module UNET_IP_maxpool_run_max_run_max_fsm (
  clk, rst, arst_n, fsm_output, main_C_1_tr0, LOOP_CH_C_0_tr0, LOOP_HEIGHT_C_0_tr0,
      LOOP_WIDTH_C_0_tr0, LOOP_Y_C_0_tr0, LOOP_X_C_0_tr0, LOOP_WIDTH_C_3_tr0, LOOP_HEIGHT_C_1_tr0,
      LOOP_CH_C_1_tr0
);
  input clk;
  input rst;
  input arst_n;
  output [12:0] fsm_output;
  reg [12:0] fsm_output;
  input main_C_1_tr0;
  input LOOP_CH_C_0_tr0;
  input LOOP_HEIGHT_C_0_tr0;
  input LOOP_WIDTH_C_0_tr0;
  input LOOP_Y_C_0_tr0;
  input LOOP_X_C_0_tr0;
  input LOOP_WIDTH_C_3_tr0;
  input LOOP_HEIGHT_C_1_tr0;
  input LOOP_CH_C_1_tr0;


  // FSM State Type Declaration for UNET_IP_maxpool_run_max_run_max_fsm_1
  parameter
    main_C_0 = 4'd0,
    main_C_1 = 4'd1,
    LOOP_CH_C_0 = 4'd2,
    LOOP_HEIGHT_C_0 = 4'd3,
    LOOP_WIDTH_C_0 = 4'd4,
    LOOP_Y_C_0 = 4'd5,
    LOOP_X_C_0 = 4'd6,
    LOOP_WIDTH_C_1 = 4'd7,
    LOOP_WIDTH_C_2 = 4'd8,
    LOOP_WIDTH_C_3 = 4'd9,
    LOOP_HEIGHT_C_1 = 4'd10,
    LOOP_CH_C_1 = 4'd11,
    main_C_2 = 4'd12;

  reg [3:0] state_var;
  reg [3:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : UNET_IP_maxpool_run_max_run_max_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 13'b0000000000010;
        if ( main_C_1_tr0 ) begin
          state_var_NS = main_C_2;
        end
        else begin
          state_var_NS = LOOP_CH_C_0;
        end
      end
      LOOP_CH_C_0 : begin
        fsm_output = 13'b0000000000100;
        if ( LOOP_CH_C_0_tr0 ) begin
          state_var_NS = LOOP_CH_C_1;
        end
        else begin
          state_var_NS = LOOP_HEIGHT_C_0;
        end
      end
      LOOP_HEIGHT_C_0 : begin
        fsm_output = 13'b0000000001000;
        if ( LOOP_HEIGHT_C_0_tr0 ) begin
          state_var_NS = LOOP_HEIGHT_C_1;
        end
        else begin
          state_var_NS = LOOP_WIDTH_C_0;
        end
      end
      LOOP_WIDTH_C_0 : begin
        fsm_output = 13'b0000000010000;
        if ( LOOP_WIDTH_C_0_tr0 ) begin
          state_var_NS = LOOP_WIDTH_C_1;
        end
        else begin
          state_var_NS = LOOP_Y_C_0;
        end
      end
      LOOP_Y_C_0 : begin
        fsm_output = 13'b0000000100000;
        if ( LOOP_Y_C_0_tr0 ) begin
          state_var_NS = LOOP_X_C_0;
        end
        else begin
          state_var_NS = LOOP_Y_C_0;
        end
      end
      LOOP_X_C_0 : begin
        fsm_output = 13'b0000001000000;
        if ( LOOP_X_C_0_tr0 ) begin
          state_var_NS = LOOP_WIDTH_C_1;
        end
        else begin
          state_var_NS = LOOP_Y_C_0;
        end
      end
      LOOP_WIDTH_C_1 : begin
        fsm_output = 13'b0000010000000;
        state_var_NS = LOOP_WIDTH_C_2;
      end
      LOOP_WIDTH_C_2 : begin
        fsm_output = 13'b0000100000000;
        state_var_NS = LOOP_WIDTH_C_3;
      end
      LOOP_WIDTH_C_3 : begin
        fsm_output = 13'b0001000000000;
        if ( LOOP_WIDTH_C_3_tr0 ) begin
          state_var_NS = LOOP_HEIGHT_C_1;
        end
        else begin
          state_var_NS = LOOP_WIDTH_C_0;
        end
      end
      LOOP_HEIGHT_C_1 : begin
        fsm_output = 13'b0010000000000;
        if ( LOOP_HEIGHT_C_1_tr0 ) begin
          state_var_NS = LOOP_CH_C_1;
        end
        else begin
          state_var_NS = LOOP_HEIGHT_C_0;
        end
      end
      LOOP_CH_C_1 : begin
        fsm_output = 13'b0100000000000;
        if ( LOOP_CH_C_1_tr0 ) begin
          state_var_NS = main_C_2;
        end
        else begin
          state_var_NS = LOOP_CH_C_0;
        end
      end
      main_C_2 : begin
        fsm_output = 13'b1000000000000;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 13'b0000000000001;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= main_C_0;
    end
    else if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    UNET_IP_maxpool_run_max
// ------------------------------------------------------------------


module UNET_IP_maxpool_run_max (
  clk, rst, arst_n, input_triosy_lz, output_triosy_lz, channels, height, width, pool_size,
      stride, input_rsci_q_d, input_rsci_radr_d, output_rsci_d_d, output_rsci_wadr_d,
      input_rsci_re_d_pff, output_rsci_we_d_pff
);
  input clk;
  input rst;
  input arst_n;
  output input_triosy_lz;
  output output_triosy_lz;
  input [6:0] channels;
  input [6:0] height;
  input [6:0] width;
  input [2:0] pool_size;
  input [2:0] stride;
  input [11:0] input_rsci_q_d;
  output [14:0] input_rsci_radr_d;
  wire [15:0] nl_input_rsci_radr_d;
  output [11:0] output_rsci_d_d;
  output [14:0] output_rsci_wadr_d;
  wire [15:0] nl_output_rsci_wadr_d;
  output input_rsci_re_d_pff;
  output output_rsci_we_d_pff;


  // Interconnect Declarations
  wire [12:0] fsm_output;
  wire and_dcpl_20;
  wire or_dcpl_21;
  reg LOOP_Y_stage_0;
  wire exit_LOOP_CH_sva_mx0;
  wire exit_LOOP_HEIGHT_sva_mx0;
  wire exit_LOOP_X_sva_mx0;
  reg [2:0] y_sva;
  reg [2:0] x_sva;
  reg exit_LOOP_Y_sva_st_2;
  reg LOOP_Y_stage_0_3;
  reg LOOP_Y_stage_0_2;
  reg exit_LOOP_Y_sva_st_1;
  reg LOOP_Y_land_lpi_6_dfm_1;
  reg LOOP_Y_stage_0_4;
  reg LOOP_Y_asn_3_itm_3;
  reg LOOP_Y_land_lpi_6_dfm_3;
  reg LOOP_Y_land_lpi_6_dfm_2;
  reg reg_input_triosy_obj_ld_cse;
  wire nor_13_cse;
  wire or_23_cse;
  reg [11:0] max_val_13_2_lpi_5;
  reg [13:0] LOOP_WIDTH_acc_6_itm;
  wire [14:0] nl_LOOP_WIDTH_acc_6_itm;
  reg [13:0] LOOP_WIDTH_mul_1_itm;
  wire [13:0] z_out_4;
  wire [14:0] z_out_5;
  wire [20:0] nl_z_out_5;
  reg [6:0] c_sva;
  reg [11:0] max_val_13_2_lpi_3;
  reg [6:0] i_sva;
  reg [6:0] j_sva;
  reg [9:0] LOOP_Y_if_acc_2_itm_1;
  wire [10:0] nl_LOOP_Y_if_acc_2_itm_1;
  reg [2:0] LOOP_Y_else_asn_itm_1;
  wire [6:0] c_sva_2;
  wire [7:0] nl_c_sva_2;
  wire [6:0] i_sva_2;
  wire [7:0] nl_i_sva_2;
  wire [6:0] j_sva_2;
  wire [7:0] nl_j_sva_2;
  wire [2:0] x_sva_2;
  wire [3:0] nl_x_sva_2;
  wire [9:0] LOOP_Y_if_mul_4_ncse_sva_1;
  reg [14:0] reg_LOOP_Y_if_acc_4_itm_1_cse;
  wire [15:0] nl_reg_LOOP_Y_if_acc_4_itm_1_cse;
  wire x_or_cse;
  wire LOOP_Y_else_if_acc_itm_12_1;
  wire LOOP_Y_acc_2_itm_3_1;
  reg z_out_6;
  reg z_out_5_1;
  reg z_out_4_1;
  reg z_out_3;
  reg z_out_2;
  reg z_out_1;
  reg z_out_0;
  reg reg_out_width_ftd;
  reg reg_out_width_ftd_1;
  reg reg_out_width_ftd_2;
  reg reg_out_width_ftd_3;
  reg reg_out_width_ftd_4;
  reg reg_out_width_ftd_5;
  reg reg_out_width_ftd_6;
  wire nand_ssc;
  reg reg_out_height_ftd;
  reg reg_out_height_ftd_1;
  reg reg_out_height_ftd_2;
  reg reg_out_height_ftd_3;
  reg reg_out_height_ftd_4;
  reg reg_out_height_ftd_5;
  reg reg_out_height_ftd_6;

  wire and_58_nl;
  wire max_val_and_nl;
  wire not_73_nl;
  wire LOOP_Y_mux_4_nl;
  wire LOOP_Y_aelse_LOOP_Y_aelse_and_nl;
  wire[7:0] LOOP_WIDTH_acc_7_nl;
  wire[8:0] nl_LOOP_WIDTH_acc_7_nl;
  wire[2:0] LOOP_Y_acc_1_nl;
  wire[3:0] nl_LOOP_Y_acc_1_nl;
  wire[14:0] LOOP_Y_if_mul_5_nl;
  wire[16:0] nl_LOOP_Y_if_mul_5_nl;
  wire[9:0] LOOP_Y_if_mux_5_nl;
  wire[9:0] LOOP_Y_else_acc_7_nl;
  wire[10:0] nl_LOOP_Y_else_acc_7_nl;
  wire and_146_nl;
  wire[6:0] LOOP_Y_if_mux_6_nl;
  wire[7:0] LOOP_CH_acc_2_nl;
  wire[8:0] nl_LOOP_CH_acc_2_nl;
  wire[7:0] LOOP_CH_acc_3_nl;
  wire[8:0] nl_LOOP_CH_acc_3_nl;
  wire[7:0] LOOP_HEIGHT_acc_2_nl;
  wire[8:0] nl_LOOP_HEIGHT_acc_2_nl;
  wire[7:0] LOOP_HEIGHT_acc_3_nl;
  wire[8:0] nl_LOOP_HEIGHT_acc_3_nl;
  wire[3:0] LOOP_X_acc_2_nl;
  wire[4:0] nl_LOOP_X_acc_2_nl;
  wire[3:0] LOOP_X_acc_3_nl;
  wire[4:0] nl_LOOP_X_acc_3_nl;
  wire[12:0] LOOP_Y_else_if_acc_nl;
  wire[3:0] LOOP_Y_acc_2_nl;
  wire[4:0] nl_LOOP_Y_acc_2_nl;
  wire[3:0] LOOP_Y_if_LOOP_Y_if_and_1_nl;
  wire[2:0] LOOP_Y_if_mux_7_nl;
  wire[6:0] LOOP_Y_if_mux_8_nl;

  // Interconnect Declarations for Component Instantiations 
  wire[7:0] LOOP_WIDTH_acc_5_nl;
  wire[8:0] nl_LOOP_WIDTH_acc_5_nl;
  wire  nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0;
  assign nl_LOOP_WIDTH_acc_5_nl = ({1'b1 , (~ reg_out_width_ftd) , (~ reg_out_width_ftd_1)
      , (~ reg_out_width_ftd_2) , (~ reg_out_width_ftd_3) , (~ reg_out_width_ftd_4)
      , (~ reg_out_width_ftd_5) , (~ reg_out_width_ftd_6)}) + 8'b00000001;
  assign LOOP_WIDTH_acc_5_nl = nl_LOOP_WIDTH_acc_5_nl[7:0];
  assign nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0 = ~ (readslicef_8_1_7(LOOP_WIDTH_acc_5_nl));
  wire  nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0;
  assign nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0 = ~(LOOP_Y_stage_0_3
      | LOOP_Y_stage_0_2 | LOOP_Y_stage_0);
  mgc_io_sync_v2 #(.valid(32'sd0)) input_triosy_obj (
      .ld(reg_input_triosy_obj_ld_cse),
      .lz(input_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) output_triosy_obj (
      .ld(reg_input_triosy_obj_ld_cse),
      .lz(output_triosy_lz)
    );
  UNET_IP_maxpool_run_max_run_max_fsm UNET_IP_maxpool_run_max_run_max_fsm_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .fsm_output(fsm_output),
      .main_C_1_tr0(exit_LOOP_CH_sva_mx0),
      .LOOP_CH_C_0_tr0(exit_LOOP_HEIGHT_sva_mx0),
      .LOOP_HEIGHT_C_0_tr0(nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0),
      .LOOP_WIDTH_C_0_tr0(exit_LOOP_X_sva_mx0),
      .LOOP_Y_C_0_tr0(nl_UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0),
      .LOOP_X_C_0_tr0(exit_LOOP_X_sva_mx0),
      .LOOP_WIDTH_C_3_tr0(LOOP_Y_stage_0),
      .LOOP_HEIGHT_C_1_tr0(exit_LOOP_HEIGHT_sva_mx0),
      .LOOP_CH_C_1_tr0(exit_LOOP_CH_sva_mx0)
    );
  assign nor_13_cse = ~(LOOP_Y_else_if_acc_itm_12_1 | LOOP_Y_land_lpi_6_dfm_3);
  assign or_23_cse = (fsm_output[1]) | (fsm_output[11]);
  assign nand_ssc = ~(and_dcpl_20 & (~ (fsm_output[1])));
  assign x_or_cse = (fsm_output[4]) | (fsm_output[6]);
  assign nl_LOOP_CH_acc_2_nl = ({1'b1 , (~ channels)}) + 8'b00000001;
  assign LOOP_CH_acc_2_nl = nl_LOOP_CH_acc_2_nl[7:0];
  assign nl_LOOP_CH_acc_3_nl = ({1'b1 , c_sva_2}) + conv_u2u_7_8(~ channels) + 8'b00000001;
  assign LOOP_CH_acc_3_nl = nl_LOOP_CH_acc_3_nl[7:0];
  assign exit_LOOP_CH_sva_mx0 = MUX_s_1_2_2((~ (readslicef_8_1_7(LOOP_CH_acc_2_nl))),
      (~ (readslicef_8_1_7(LOOP_CH_acc_3_nl))), fsm_output[11]);
  assign nl_c_sva_2 = c_sva + 7'b0000001;
  assign c_sva_2 = nl_c_sva_2[6:0];
  assign nl_LOOP_HEIGHT_acc_2_nl = ({1'b1 , (~ reg_out_height_ftd) , (~ reg_out_height_ftd_1)
      , (~ reg_out_height_ftd_2) , (~ reg_out_height_ftd_3) , (~ reg_out_height_ftd_4)
      , (~ reg_out_height_ftd_5) , (~ reg_out_height_ftd_6)}) + 8'b00000001;
  assign LOOP_HEIGHT_acc_2_nl = nl_LOOP_HEIGHT_acc_2_nl[7:0];
  assign nl_LOOP_HEIGHT_acc_3_nl = ({1'b1 , i_sva_2}) + conv_u2u_7_8({(~ reg_out_height_ftd)
      , (~ reg_out_height_ftd_1) , (~ reg_out_height_ftd_2) , (~ reg_out_height_ftd_3)
      , (~ reg_out_height_ftd_4) , (~ reg_out_height_ftd_5) , (~ reg_out_height_ftd_6)})
      + 8'b00000001;
  assign LOOP_HEIGHT_acc_3_nl = nl_LOOP_HEIGHT_acc_3_nl[7:0];
  assign exit_LOOP_HEIGHT_sva_mx0 = MUX_s_1_2_2((~ (readslicef_8_1_7(LOOP_HEIGHT_acc_2_nl))),
      (~ (readslicef_8_1_7(LOOP_HEIGHT_acc_3_nl))), fsm_output[10]);
  assign nl_i_sva_2 = i_sva + 7'b0000001;
  assign i_sva_2 = nl_i_sva_2[6:0];
  assign nl_j_sva_2 = j_sva + 7'b0000001;
  assign j_sva_2 = nl_j_sva_2[6:0];
  assign nl_LOOP_X_acc_2_nl = ({1'b1 , (~ pool_size)}) + 4'b0001;
  assign LOOP_X_acc_2_nl = nl_LOOP_X_acc_2_nl[3:0];
  assign nl_LOOP_X_acc_3_nl = ({1'b1 , x_sva_2}) + conv_u2u_3_4(~ pool_size) + 4'b0001;
  assign LOOP_X_acc_3_nl = nl_LOOP_X_acc_3_nl[3:0];
  assign exit_LOOP_X_sva_mx0 = MUX_s_1_2_2((~ (readslicef_4_1_3(LOOP_X_acc_2_nl))),
      (~ (readslicef_4_1_3(LOOP_X_acc_3_nl))), fsm_output[6]);
  assign nl_x_sva_2 = x_sva + 3'b001;
  assign x_sva_2 = nl_x_sva_2[2:0];
  assign LOOP_Y_if_mul_4_ncse_sva_1 = j_sva * stride;
  assign LOOP_Y_else_if_acc_nl = $signed(max_val_13_2_lpi_3) - $signed(input_rsci_q_d);
  assign LOOP_Y_else_if_acc_itm_12_1 = readslicef_13_1_12(LOOP_Y_else_if_acc_nl);
  assign and_dcpl_20 = ~((fsm_output[0]) | (fsm_output[12]));
  assign or_dcpl_21 = (fsm_output[9]) | (fsm_output[6]) | (fsm_output[8]);
  assign nl_LOOP_Y_acc_2_nl = ({1'b1 , y_sva}) + conv_u2u_3_4(~ pool_size) + 4'b0001;
  assign LOOP_Y_acc_2_nl = nl_LOOP_Y_acc_2_nl[3:0];
  assign LOOP_Y_acc_2_itm_3_1 = readslicef_4_1_3(LOOP_Y_acc_2_nl);
  assign nl_input_rsci_radr_d = reg_LOOP_Y_if_acc_4_itm_1_cse + z_out_5;
  assign input_rsci_radr_d = nl_input_rsci_radr_d[14:0];
  assign input_rsci_re_d_pff = (~ exit_LOOP_Y_sva_st_2) & LOOP_Y_stage_0_3 & (fsm_output[5]);
  assign output_rsci_d_d = max_val_13_2_lpi_5;
  assign nl_output_rsci_wadr_d = conv_u2u_14_15(LOOP_WIDTH_acc_6_itm) + z_out_5;
  assign output_rsci_wadr_d = nl_output_rsci_wadr_d[14:0];
  assign output_rsci_we_d_pff = fsm_output[8];
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd <= z_out_6;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_1 <= z_out_5_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_2 <= z_out_4_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_3 <= z_out_3;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_4 <= z_out_2;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_5 <= z_out_1;
    end
  end
  always @(posedge clk) begin
    if ( ~ and_dcpl_20 ) begin
      reg_out_width_ftd_6 <= z_out_0;
    end
  end
  always @(posedge clk) begin
    if ( (~(((fsm_output[9:5]==5'b00000)) | ((nor_13_cse | LOOP_Y_asn_3_itm_3 | (~
        LOOP_Y_stage_0_4)) & (fsm_output[5])))) | (fsm_output[4]) ) begin
      max_val_13_2_lpi_3 <= MUX_v_12_2_2(max_val_13_2_lpi_5, input_rsci_q_d, and_58_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_input_triosy_obj_ld_cse <= 1'b0;
      LOOP_Y_asn_3_itm_3 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_3 <= 1'b0;
      exit_LOOP_Y_sva_st_2 <= 1'b0;
      exit_LOOP_Y_sva_st_1 <= 1'b0;
      y_sva <= 3'b000;
      LOOP_Y_stage_0_2 <= 1'b0;
      LOOP_Y_stage_0_3 <= 1'b0;
      LOOP_Y_stage_0_4 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_2 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_1 <= 1'b0;
    end
    else if ( rst ) begin
      reg_input_triosy_obj_ld_cse <= 1'b0;
      LOOP_Y_asn_3_itm_3 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_3 <= 1'b0;
      exit_LOOP_Y_sva_st_2 <= 1'b0;
      exit_LOOP_Y_sva_st_1 <= 1'b0;
      y_sva <= 3'b000;
      LOOP_Y_stage_0_2 <= 1'b0;
      LOOP_Y_stage_0_3 <= 1'b0;
      LOOP_Y_stage_0_4 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_2 <= 1'b0;
      LOOP_Y_land_lpi_6_dfm_1 <= 1'b0;
    end
    else begin
      reg_input_triosy_obj_ld_cse <= exit_LOOP_CH_sva_mx0 & or_23_cse;
      LOOP_Y_asn_3_itm_3 <= exit_LOOP_Y_sva_st_2;
      LOOP_Y_land_lpi_6_dfm_3 <= LOOP_Y_land_lpi_6_dfm_2;
      exit_LOOP_Y_sva_st_2 <= exit_LOOP_Y_sva_st_1;
      exit_LOOP_Y_sva_st_1 <= ~ LOOP_Y_acc_2_itm_3_1;
      y_sva <= MUX_v_3_2_2(3'b000, LOOP_Y_acc_1_nl, (fsm_output[5]));
      LOOP_Y_stage_0_2 <= LOOP_Y_stage_0 & (fsm_output[5]);
      LOOP_Y_stage_0_3 <= LOOP_Y_stage_0_2 & (fsm_output[5]);
      LOOP_Y_stage_0_4 <= LOOP_Y_stage_0_3 & (fsm_output[5]);
      LOOP_Y_land_lpi_6_dfm_2 <= LOOP_Y_land_lpi_6_dfm_1;
      LOOP_Y_land_lpi_6_dfm_1 <= ~((y_sva!=3'b000) | (x_sva!=3'b000));
    end
  end
  always @(posedge clk) begin
    if ( or_23_cse ) begin
      c_sva <= MUX_v_7_2_2(7'b0000000, c_sva_2, (fsm_output[11]));
    end
  end
  always @(posedge clk) begin
    if ( nand_ssc ) begin
      reg_out_height_ftd <= z_out_6;
      reg_out_height_ftd_1 <= z_out_5_1;
      reg_out_height_ftd_2 <= z_out_4_1;
      reg_out_height_ftd_3 <= z_out_3;
      reg_out_height_ftd_4 <= z_out_2;
      reg_out_height_ftd_5 <= z_out_1;
      reg_out_height_ftd_6 <= z_out_0;
    end
  end
  always @(posedge clk) begin
    if ( (fsm_output[10]) | (fsm_output[2]) ) begin
      i_sva <= MUX_v_7_2_2(7'b0000000, i_sva_2, (fsm_output[10]));
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_21 | (fsm_output[4]) | (fsm_output[7])) ) begin
      max_val_13_2_lpi_5 <= MUX_v_12_2_2(max_val_13_2_lpi_3, input_rsci_q_d, max_val_and_nl);
    end
  end
  always @(posedge clk) begin
    if ( ~(or_dcpl_21 | (fsm_output[5:4]!=2'b00)) ) begin
      j_sva <= MUX_v_7_2_2(7'b0000000, j_sva_2, not_73_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      x_sva <= 3'b000;
    end
    else if ( rst ) begin
      x_sva <= 3'b000;
    end
    else if ( x_or_cse ) begin
      x_sva <= MUX_v_3_2_2(3'b000, x_sva_2, (fsm_output[6]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      LOOP_Y_stage_0 <= 1'b0;
    end
    else if ( rst ) begin
      LOOP_Y_stage_0 <= 1'b0;
    end
    else if ( x_or_cse | (fsm_output[5]) | (fsm_output[7]) ) begin
      LOOP_Y_stage_0 <= LOOP_Y_mux_4_nl | x_or_cse;
    end
  end
  always @(posedge clk) begin
    reg_LOOP_Y_if_acc_4_itm_1_cse <= nl_reg_LOOP_Y_if_acc_4_itm_1_cse[14:0];
    LOOP_Y_else_asn_itm_1 <= y_sva;
    LOOP_Y_if_acc_2_itm_1 <= nl_LOOP_Y_if_acc_2_itm_1[9:0];
    LOOP_WIDTH_mul_1_itm <= c_sva * LOOP_Y_if_mux_6_nl;
    LOOP_WIDTH_acc_6_itm <= nl_LOOP_WIDTH_acc_6_itm[13:0];
  end
  assign and_58_nl = (LOOP_Y_else_if_acc_itm_12_1 | LOOP_Y_land_lpi_6_dfm_3) & (~
      LOOP_Y_asn_3_itm_3) & LOOP_Y_stage_0_4 & (fsm_output[5]);
  assign nl_LOOP_Y_acc_1_nl = y_sva + 3'b001;
  assign LOOP_Y_acc_1_nl = nl_LOOP_Y_acc_1_nl[2:0];
  assign max_val_and_nl = (~((nor_13_cse | LOOP_Y_asn_3_itm_3) & LOOP_Y_stage_0_4))
      & (fsm_output[5]);
  assign not_73_nl = ~ (fsm_output[3]);
  assign LOOP_Y_aelse_LOOP_Y_aelse_and_nl = LOOP_Y_stage_0 & LOOP_Y_acc_2_itm_3_1;
  assign nl_LOOP_WIDTH_acc_7_nl = ({1'b1 , j_sva_2}) + conv_u2u_7_8({(~ reg_out_width_ftd)
      , (~ reg_out_width_ftd_1) , (~ reg_out_width_ftd_2) , (~ reg_out_width_ftd_3)
      , (~ reg_out_width_ftd_4) , (~ reg_out_width_ftd_5) , (~ reg_out_width_ftd_6)})
      + 8'b00000001;
  assign LOOP_WIDTH_acc_7_nl = nl_LOOP_WIDTH_acc_7_nl[7:0];
  assign LOOP_Y_mux_4_nl = MUX_s_1_2_2(LOOP_Y_aelse_LOOP_Y_aelse_and_nl, (~ (readslicef_8_1_7(LOOP_WIDTH_acc_7_nl))),
      fsm_output[7]);
  assign nl_LOOP_Y_if_mul_5_nl = LOOP_Y_if_acc_2_itm_1 * width;
  assign LOOP_Y_if_mul_5_nl = nl_LOOP_Y_if_mul_5_nl[14:0];
  assign nl_LOOP_Y_else_acc_7_nl = LOOP_Y_if_mul_4_ncse_sva_1 + conv_u2u_3_10(LOOP_Y_else_asn_itm_1);
  assign LOOP_Y_else_acc_7_nl = nl_LOOP_Y_else_acc_7_nl[9:0];
  assign and_146_nl = (~ LOOP_Y_land_lpi_6_dfm_1) & (fsm_output[5]);
  assign LOOP_Y_if_mux_5_nl = MUX_v_10_2_2(LOOP_Y_if_mul_4_ncse_sva_1, LOOP_Y_else_acc_7_nl,
      and_146_nl);
  assign nl_reg_LOOP_Y_if_acc_4_itm_1_cse  = LOOP_Y_if_mul_5_nl + conv_u2u_10_15(LOOP_Y_if_mux_5_nl);
  assign nl_LOOP_Y_if_acc_2_itm_1  = (z_out_4[9:0]) + conv_u2u_3_10(x_sva);
  assign LOOP_Y_if_mux_6_nl = MUX_v_7_2_2(height, ({reg_out_height_ftd , reg_out_height_ftd_1
      , reg_out_height_ftd_2 , reg_out_height_ftd_3 , reg_out_height_ftd_4 , reg_out_height_ftd_5
      , reg_out_height_ftd_6}), fsm_output[7]);
  assign nl_LOOP_WIDTH_acc_6_itm  = z_out_4 + conv_u2u_7_14(j_sva);
  always @(width or height or fsm_output or stride)
  begin : mgc_div_7_3_0_b0_line_26
    // Interconnect Declarations
    reg [3:0] divmod6448_2_diff_1;
    reg [3:0] divmod6448_2_diff_2;
    reg [3:0] divmod6448_2_diff_3;
    reg [3:0] divmod6448_2_diff_4;
    reg [3:0] divmod6448_2_diff_5;
    reg [3:0] divmod6448_2_diff_6;
    reg divmod6448_2_lbuf_8_3;
    reg divmod6448_2_lbuf_8_4;
    reg divmod6448_2_lbuf_8_5;
    reg divmod6448_2_lbuf_8_6;
    reg divmod6448_2_lbuf_7_2;
    reg divmod6448_2_lbuf_7_3;
    reg divmod6448_2_lbuf_7_4;
    reg divmod6448_2_lbuf_7_5;
    reg divmod6448_2_lbuf_7_6;
    reg divmod6448_2_lbuf_6;
    reg divmod6448_2_lbuf_6_1;
    reg divmod6448_2_lbuf_6_2;
    reg divmod6448_2_lbuf_6_3;
    reg divmod6448_2_lbuf_6_4;
    reg slc_fsm_output_1_5_ssc;
    reg divmod6448_2_lbuf_6_5;
    reg [5:0] divmod6448_2_lbuf_5_0;

    reg[3:0] divmod6448_2_loop951_7_acc_1_nl;
    reg[5:0] nl_divmod6448_2_loop951_7_acc_1_nl;
    slc_fsm_output_1_5_ssc = fsm_output[1];
    divmod6448_2_lbuf_5_0 = MUX_v_6_2_2((width[5:0]), (height[5:0]), slc_fsm_output_1_5_ssc);
    divmod6448_2_lbuf_6_5 = MUX_s_1_2_2((width[6]), (height[6]), slc_fsm_output_1_5_ssc);
    divmod6448_2_diff_1 = conv_u2u_1_4(divmod6448_2_lbuf_6_5) + ({1'b1 , (~ stride)})
        + 4'b0001;
    if ( divmod6448_2_diff_1[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_6_5 = divmod6448_2_diff_1[0];
    end
    divmod6448_2_lbuf_7_2 = divmod6448_2_lbuf_6_5;
    divmod6448_2_lbuf_6 = divmod6448_2_lbuf_5_0[5];
    divmod6448_2_diff_2 = conv_u2u_2_4({divmod6448_2_lbuf_6_5 , (divmod6448_2_lbuf_5_0[5])})
        + ({1'b1 , (~ stride)}) + 4'b0001;
    if ( divmod6448_2_diff_2[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_7_2 = divmod6448_2_diff_2[1];
      divmod6448_2_lbuf_6 = divmod6448_2_diff_2[0];
    end
    divmod6448_2_lbuf_8_3 = divmod6448_2_lbuf_7_2;
    divmod6448_2_lbuf_7_3 = divmod6448_2_lbuf_6;
    divmod6448_2_lbuf_6_1 = divmod6448_2_lbuf_5_0[4];
    divmod6448_2_diff_3 = conv_u2u_3_4({divmod6448_2_lbuf_7_2 , divmod6448_2_lbuf_6
        , (divmod6448_2_lbuf_5_0[4])}) + ({1'b1 , (~ stride)}) + 4'b0001;
    if ( divmod6448_2_diff_3[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_7_3 = divmod6448_2_diff_3[1];
      divmod6448_2_lbuf_8_3 = divmod6448_2_diff_3[2];
      divmod6448_2_lbuf_6_1 = divmod6448_2_diff_3[0];
    end
    divmod6448_2_lbuf_8_4 = divmod6448_2_lbuf_7_3;
    divmod6448_2_lbuf_7_4 = divmod6448_2_lbuf_6_1;
    divmod6448_2_lbuf_6_2 = divmod6448_2_lbuf_5_0[3];
    divmod6448_2_diff_4 = ({divmod6448_2_lbuf_8_3 , divmod6448_2_lbuf_7_3 , divmod6448_2_lbuf_6_1
        , (divmod6448_2_lbuf_5_0[3])}) + ({1'b1 , (~ stride)}) + 4'b0001;
    if ( divmod6448_2_diff_4[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_7_4 = divmod6448_2_diff_4[1];
      divmod6448_2_lbuf_8_4 = divmod6448_2_diff_4[2];
      divmod6448_2_lbuf_6_2 = divmod6448_2_diff_4[0];
    end
    divmod6448_2_lbuf_8_5 = divmod6448_2_lbuf_7_4;
    divmod6448_2_lbuf_7_5 = divmod6448_2_lbuf_6_2;
    divmod6448_2_lbuf_6_3 = divmod6448_2_lbuf_5_0[2];
    divmod6448_2_diff_5 = ({divmod6448_2_lbuf_8_4 , divmod6448_2_lbuf_7_4 , divmod6448_2_lbuf_6_2
        , (divmod6448_2_lbuf_5_0[2])}) + ({1'b1 , (~ stride)}) + 4'b0001;
    if ( divmod6448_2_diff_5[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_7_5 = divmod6448_2_diff_5[1];
      divmod6448_2_lbuf_8_5 = divmod6448_2_diff_5[2];
      divmod6448_2_lbuf_6_3 = divmod6448_2_diff_5[0];
    end
    divmod6448_2_lbuf_8_6 = divmod6448_2_lbuf_7_5;
    divmod6448_2_lbuf_7_6 = divmod6448_2_lbuf_6_3;
    divmod6448_2_lbuf_6_4 = divmod6448_2_lbuf_5_0[1];
    divmod6448_2_diff_6 = ({divmod6448_2_lbuf_8_5 , divmod6448_2_lbuf_7_5 , divmod6448_2_lbuf_6_3
        , (divmod6448_2_lbuf_5_0[1])}) + ({1'b1 , (~ stride)}) + 4'b0001;
    if ( divmod6448_2_diff_6[3] ) begin
    end
    else begin
      divmod6448_2_lbuf_7_6 = divmod6448_2_diff_6[1];
      divmod6448_2_lbuf_8_6 = divmod6448_2_diff_6[2];
      divmod6448_2_lbuf_6_4 = divmod6448_2_diff_6[0];
    end
    z_out_3 = ~ (divmod6448_2_diff_4[3]);
    z_out_2 = ~ (divmod6448_2_diff_5[3]);
    z_out_4_1 = ~ (divmod6448_2_diff_3[3]);
    z_out_1 = ~ (divmod6448_2_diff_6[3]);
    z_out_5_1 = ~ (divmod6448_2_diff_2[3]);
    nl_divmod6448_2_loop951_7_acc_1_nl = ({divmod6448_2_lbuf_8_6 , divmod6448_2_lbuf_7_6
        , divmod6448_2_lbuf_6_4 , (divmod6448_2_lbuf_5_0[0])}) + ({1'b1 , (~ stride)})
        + 4'b0001;
    divmod6448_2_loop951_7_acc_1_nl = nl_divmod6448_2_loop951_7_acc_1_nl[3:0];
    z_out_0 = ~ (readslicef_4_1_3(divmod6448_2_loop951_7_acc_1_nl));
    z_out_6 = ~ (divmod6448_2_diff_1[3]);
  end

  assign LOOP_Y_if_LOOP_Y_if_and_1_nl = MUX_v_4_2_2(4'b0000, ({reg_out_width_ftd
      , reg_out_width_ftd_1 , reg_out_width_ftd_2 , reg_out_width_ftd_3}), (fsm_output[7]));
  assign LOOP_Y_if_mux_7_nl = MUX_v_3_2_2(stride, ({reg_out_width_ftd_4 , reg_out_width_ftd_5
      , reg_out_width_ftd_6}), fsm_output[7]);
  assign z_out_4 = i_sva * ({LOOP_Y_if_LOOP_Y_if_and_1_nl , LOOP_Y_if_mux_7_nl});
  assign LOOP_Y_if_mux_8_nl = MUX_v_7_2_2(width, ({reg_out_width_ftd , reg_out_width_ftd_1
      , reg_out_width_ftd_2 , reg_out_width_ftd_3 , reg_out_width_ftd_4 , reg_out_width_ftd_5
      , reg_out_width_ftd_6}), fsm_output[8]);
  assign nl_z_out_5 = LOOP_Y_if_mux_8_nl * LOOP_WIDTH_mul_1_itm;
  assign z_out_5 = nl_z_out_5[14:0];

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [9:0] MUX_v_10_2_2;
    input [9:0] input_0;
    input [9:0] input_1;
    input  sel;
    reg [9:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_10_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_13_1_12;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 12;
    readslicef_13_1_12 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [3:0] conv_u2u_1_4 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_4 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [9:0] conv_u2u_3_10 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_10 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction


  function automatic [13:0] conv_u2u_7_14 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_14 = {{7{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_10_15 ;
    input [9:0]  vector ;
  begin
    conv_u2u_10_15 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [14:0] conv_u2u_14_15 ;
    input [13:0]  vector ;
  begin
    conv_u2u_14_15 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    UNET_IP_maxpool
// ------------------------------------------------------------------


module UNET_IP_maxpool (
  clk, rst, arst_n, input_rsc_radr, input_rsc_re, input_rsc_q, input_rsc_clken, input_triosy_lz,
      output_rsc_wadr, output_rsc_d, output_rsc_we, output_rsc_clken, output_triosy_lz,
      channels, height, width, pool_size, stride
);
  input clk;
  input rst;
  input arst_n;
  output [14:0] input_rsc_radr;
  output input_rsc_re;
  input [11:0] input_rsc_q;
  output input_rsc_clken;
  output input_triosy_lz;
  output [14:0] output_rsc_wadr;
  output [11:0] output_rsc_d;
  output output_rsc_we;
  output output_rsc_clken;
  output output_triosy_lz;
  input [6:0] channels;
  input [6:0] height;
  input [6:0] width;
  input [2:0] pool_size;
  input [2:0] stride;


  // Interconnect Declarations
  wire [11:0] input_rsci_q_d;
  wire [14:0] input_rsci_radr_d;
  wire [11:0] output_rsci_d_d;
  wire [14:0] output_rsci_wadr_d;
  wire input_rsci_re_d_iff;
  wire output_rsci_we_d_iff;


  // Interconnect Declarations for Component Instantiations 
  UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
      input_rsci (
      .clken(input_rsc_clken),
      .q(input_rsc_q),
      .re(input_rsc_re),
      .radr(input_rsc_radr),
      .clken_d(1'b1),
      .q_d(input_rsci_q_d),
      .radr_d(input_rsci_radr_d),
      .re_d(input_rsci_re_d_iff),
      .readA_r_ram_ir_internal_RMASK_B_d(input_rsci_re_d_iff)
    );
  UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
      output_rsci (
      .clken(output_rsc_clken),
      .we(output_rsc_we),
      .d(output_rsc_d),
      .wadr(output_rsc_wadr),
      .clken_d(1'b1),
      .d_d(output_rsci_d_d),
      .wadr_d(output_rsci_wadr_d),
      .we_d(output_rsci_we_d_iff),
      .writeA_w_ram_ir_internal_WMASK_B_d(output_rsci_we_d_iff)
    );
  UNET_IP_maxpool_run_max UNET_IP_maxpool_run_max_inst (
      .clk(clk),
      .rst(rst),
      .arst_n(arst_n),
      .input_triosy_lz(input_triosy_lz),
      .output_triosy_lz(output_triosy_lz),
      .channels(channels),
      .height(height),
      .width(width),
      .pool_size(pool_size),
      .stride(stride),
      .input_rsci_q_d(input_rsci_q_d),
      .input_rsci_radr_d(input_rsci_radr_d),
      .output_rsci_d_d(output_rsci_d_d),
      .output_rsci_wadr_d(output_rsci_wadr_d),
      .input_rsci_re_d_pff(input_rsci_re_d_iff),
      .output_rsci_we_d_pff(output_rsci_we_d_iff)
    );
endmodule



