
--------> /home/raid7_4/raid1_1/linux/mentor/Catapult/2023.2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.vhd 
--------------------------------------------------------------------------------
-- Catapult Synthesis - Sample I/O Port Library
--
-- Copyright (c) 2003-2017 Mentor Graphics Corp.
--       All Rights Reserved
--
-- This document may be used and distributed without restriction provided that
-- this copyright statement is not removed from the file and that any derivative
-- work contains this copyright notice.
--
-- The design information contained in this file is intended to be an example
-- of the functionality which the end user may study in preparation for creating
-- their own custom interfaces. This design does not necessarily present a 
-- complete implementation of the named protocol or standard.
--
--------------------------------------------------------------------------------

LIBRARY ieee;

USE ieee.std_logic_1164.all;
PACKAGE mgc_io_sync_pkg_v2 IS

COMPONENT mgc_io_sync_v2
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END COMPONENT;

END mgc_io_sync_pkg_v2;

LIBRARY ieee;

USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all; -- Prevent STARC 2.1.1.2 violation

ENTITY mgc_io_sync_v2 IS
  GENERIC (
    valid    : INTEGER RANGE 0 TO 1
  );
  PORT (
    ld       : IN    std_logic;
    lz       : OUT   std_logic
  );
END mgc_io_sync_v2;

ARCHITECTURE beh OF mgc_io_sync_v2 IS
BEGIN

  lz <= ld;

END beh;


--------> ./rtl.vhdl 
-- ----------------------------------------------------------------------
--  HLS HDL:        VHDL Netlister
--  HLS Version:    2023.2/1059873 Production Release
--  HLS Date:       Mon Aug  7 10:54:31 PDT 2023
-- 
--  Generated by:   r12016@cad40
--  Generated date: Thu Jun 13 02:36:30 2024
-- ----------------------------------------------------------------------

-- 
-- ------------------------------------------------------------------
--  Design Unit:    UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
    IS
  PORT(
    clken : OUT STD_LOGIC;
    we : OUT STD_LOGIC;
    d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    wadr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    d_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    wadr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
    we_d : IN STD_LOGIC;
    writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
  );
END UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen;

ARCHITECTURE v1 OF UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  we <= (writeA_w_ram_ir_internal_WMASK_B_d);
  d <= (d_d);
  wadr <= (wadr_d);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
    IS
  PORT(
    clken : OUT STD_LOGIC;
    q : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    re : OUT STD_LOGIC;
    radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    clken_d : IN STD_LOGIC;
    q_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    radr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
    re_d : IN STD_LOGIC;
    readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
  );
END UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen;

ARCHITECTURE v1 OF UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
    IS
  -- Default Constants

BEGIN
  clken <= (clken_d);
  q_d <= q;
  re <= (readA_r_ram_ir_internal_RMASK_B_d);
  radr <= (radr_d);
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    UNET_IP_maxpool_run_max_run_max_fsm
--  FSM Module
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY UNET_IP_maxpool_run_max_run_max_fsm IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    arst_n : IN STD_LOGIC;
    fsm_output : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
    main_C_1_tr0 : IN STD_LOGIC;
    LOOP_CH_C_0_tr0 : IN STD_LOGIC;
    LOOP_HEIGHT_C_0_tr0 : IN STD_LOGIC;
    LOOP_WIDTH_C_0_tr0 : IN STD_LOGIC;
    LOOP_Y_C_0_tr0 : IN STD_LOGIC;
    LOOP_X_C_0_tr0 : IN STD_LOGIC;
    LOOP_WIDTH_C_3_tr0 : IN STD_LOGIC;
    LOOP_HEIGHT_C_1_tr0 : IN STD_LOGIC;
    LOOP_CH_C_1_tr0 : IN STD_LOGIC
  );
END UNET_IP_maxpool_run_max_run_max_fsm;

ARCHITECTURE v1 OF UNET_IP_maxpool_run_max_run_max_fsm IS
  -- Default Constants

  -- FSM State Type Declaration for UNET_IP_maxpool_run_max_run_max_fsm_1
  TYPE UNET_IP_maxpool_run_max_run_max_fsm_1_ST IS (main_C_0, main_C_1, LOOP_CH_C_0,
      LOOP_HEIGHT_C_0, LOOP_WIDTH_C_0, LOOP_Y_C_0, LOOP_X_C_0, LOOP_WIDTH_C_1, LOOP_WIDTH_C_2,
      LOOP_WIDTH_C_3, LOOP_HEIGHT_C_1, LOOP_CH_C_1, main_C_2);

  SIGNAL state_var : UNET_IP_maxpool_run_max_run_max_fsm_1_ST;
  SIGNAL state_var_NS : UNET_IP_maxpool_run_max_run_max_fsm_1_ST;

BEGIN
  UNET_IP_maxpool_run_max_run_max_fsm_1 : PROCESS (main_C_1_tr0, LOOP_CH_C_0_tr0,
      LOOP_HEIGHT_C_0_tr0, LOOP_WIDTH_C_0_tr0, LOOP_Y_C_0_tr0, LOOP_X_C_0_tr0, LOOP_WIDTH_C_3_tr0,
      LOOP_HEIGHT_C_1_tr0, LOOP_CH_C_1_tr0, state_var)
  BEGIN
    CASE state_var IS
      WHEN main_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000010");
        IF ( main_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_2;
        ELSE
          state_var_NS <= LOOP_CH_C_0;
        END IF;
      WHEN LOOP_CH_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000100");
        IF ( LOOP_CH_C_0_tr0 = '1' ) THEN
          state_var_NS <= LOOP_CH_C_1;
        ELSE
          state_var_NS <= LOOP_HEIGHT_C_0;
        END IF;
      WHEN LOOP_HEIGHT_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000001000");
        IF ( LOOP_HEIGHT_C_0_tr0 = '1' ) THEN
          state_var_NS <= LOOP_HEIGHT_C_1;
        ELSE
          state_var_NS <= LOOP_WIDTH_C_0;
        END IF;
      WHEN LOOP_WIDTH_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000010000");
        IF ( LOOP_WIDTH_C_0_tr0 = '1' ) THEN
          state_var_NS <= LOOP_WIDTH_C_1;
        ELSE
          state_var_NS <= LOOP_Y_C_0;
        END IF;
      WHEN LOOP_Y_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000100000");
        IF ( LOOP_Y_C_0_tr0 = '1' ) THEN
          state_var_NS <= LOOP_X_C_0;
        ELSE
          state_var_NS <= LOOP_Y_C_0;
        END IF;
      WHEN LOOP_X_C_0 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000001000000");
        IF ( LOOP_X_C_0_tr0 = '1' ) THEN
          state_var_NS <= LOOP_WIDTH_C_1;
        ELSE
          state_var_NS <= LOOP_Y_C_0;
        END IF;
      WHEN LOOP_WIDTH_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000010000000");
        state_var_NS <= LOOP_WIDTH_C_2;
      WHEN LOOP_WIDTH_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000100000000");
        state_var_NS <= LOOP_WIDTH_C_3;
      WHEN LOOP_WIDTH_C_3 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0001000000000");
        IF ( LOOP_WIDTH_C_3_tr0 = '1' ) THEN
          state_var_NS <= LOOP_HEIGHT_C_1;
        ELSE
          state_var_NS <= LOOP_WIDTH_C_0;
        END IF;
      WHEN LOOP_HEIGHT_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0010000000000");
        IF ( LOOP_HEIGHT_C_1_tr0 = '1' ) THEN
          state_var_NS <= LOOP_CH_C_1;
        ELSE
          state_var_NS <= LOOP_HEIGHT_C_0;
        END IF;
      WHEN LOOP_CH_C_1 =>
        fsm_output <= STD_LOGIC_VECTOR'( "0100000000000");
        IF ( LOOP_CH_C_1_tr0 = '1' ) THEN
          state_var_NS <= main_C_2;
        ELSE
          state_var_NS <= LOOP_CH_C_0;
        END IF;
      WHEN main_C_2 =>
        fsm_output <= STD_LOGIC_VECTOR'( "1000000000000");
        state_var_NS <= main_C_0;
      -- main_C_0
      WHEN OTHERS =>
        fsm_output <= STD_LOGIC_VECTOR'( "0000000000001");
        state_var_NS <= main_C_1;
    END CASE;
  END PROCESS UNET_IP_maxpool_run_max_run_max_fsm_1;

  UNET_IP_maxpool_run_max_run_max_fsm_1_REG : PROCESS (clk, arst_n)
  BEGIN
    IF ( arst_n = '0' ) THEN
      state_var <= main_C_0;
    ELSIF clk'event AND ( clk = '1' ) THEN
      IF ( rst = '1' ) THEN
        state_var <= main_C_0;
      ELSE
        state_var <= state_var_NS;
      END IF;
    END IF;
  END PROCESS UNET_IP_maxpool_run_max_run_max_fsm_1_REG;

END v1;

-- ------------------------------------------------------------------
--  Design Unit:    UNET_IP_maxpool_run_max
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY UNET_IP_maxpool_run_max IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    arst_n : IN STD_LOGIC;
    input_triosy_lz : OUT STD_LOGIC;
    output_triosy_lz : OUT STD_LOGIC;
    channels : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    height : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    width : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    pool_size : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    stride : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    input_rsci_q_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    input_rsci_radr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    output_rsci_d_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    output_rsci_wadr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    input_rsci_re_d_pff : OUT STD_LOGIC;
    output_rsci_we_d_pff : OUT STD_LOGIC
  );
END UNET_IP_maxpool_run_max;

ARCHITECTURE v1 OF UNET_IP_maxpool_run_max IS
  -- Default Constants

  -- Interconnect Declarations
  SIGNAL fsm_output : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL and_dcpl_20 : STD_LOGIC;
  SIGNAL or_dcpl_21 : STD_LOGIC;
  SIGNAL LOOP_Y_stage_0 : STD_LOGIC;
  SIGNAL exit_LOOP_CH_sva_mx0 : STD_LOGIC;
  SIGNAL exit_LOOP_HEIGHT_sva_mx0 : STD_LOGIC;
  SIGNAL exit_LOOP_X_sva_mx0 : STD_LOGIC;
  SIGNAL y_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL x_sva : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL exit_LOOP_Y_sva_st_2 : STD_LOGIC;
  SIGNAL LOOP_Y_stage_0_3 : STD_LOGIC;
  SIGNAL LOOP_Y_stage_0_2 : STD_LOGIC;
  SIGNAL exit_LOOP_Y_sva_st_1 : STD_LOGIC;
  SIGNAL LOOP_Y_land_lpi_6_dfm_1 : STD_LOGIC;
  SIGNAL LOOP_Y_stage_0_4 : STD_LOGIC;
  SIGNAL LOOP_Y_asn_3_itm_3 : STD_LOGIC;
  SIGNAL LOOP_Y_land_lpi_6_dfm_3 : STD_LOGIC;
  SIGNAL LOOP_Y_land_lpi_6_dfm_2 : STD_LOGIC;
  SIGNAL reg_input_triosy_obj_ld_cse : STD_LOGIC;
  SIGNAL nor_13_cse : STD_LOGIC;
  SIGNAL or_23_cse : STD_LOGIC;
  SIGNAL max_val_13_2_lpi_5 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL LOOP_WIDTH_acc_6_itm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL LOOP_WIDTH_mul_1_itm : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL z_out_4 : STD_LOGIC_VECTOR (13 DOWNTO 0);
  SIGNAL z_out_5 : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL c_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL max_val_13_2_lpi_3 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL i_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL j_sva : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL LOOP_Y_if_acc_2_itm_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL LOOP_Y_else_asn_itm_1 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL c_sva_2 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL i_sva_2 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL j_sva_2 : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL x_sva_2 : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL LOOP_Y_if_mul_4_ncse_sva_1 : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL reg_LOOP_Y_if_acc_4_itm_1_cse : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL x_or_cse : STD_LOGIC;
  SIGNAL LOOP_Y_else_if_acc_itm_12_1 : STD_LOGIC;
  SIGNAL LOOP_Y_acc_2_itm_3_1 : STD_LOGIC;
  SIGNAL z_out_6 : STD_LOGIC;
  SIGNAL z_out_5_1 : STD_LOGIC;
  SIGNAL z_out_4_1 : STD_LOGIC;
  SIGNAL z_out_3 : STD_LOGIC;
  SIGNAL z_out_2 : STD_LOGIC;
  SIGNAL z_out_1 : STD_LOGIC;
  SIGNAL z_out_0 : STD_LOGIC;
  SIGNAL reg_out_width_ftd : STD_LOGIC;
  SIGNAL reg_out_width_ftd_1 : STD_LOGIC;
  SIGNAL reg_out_width_ftd_2 : STD_LOGIC;
  SIGNAL reg_out_width_ftd_3 : STD_LOGIC;
  SIGNAL reg_out_width_ftd_4 : STD_LOGIC;
  SIGNAL reg_out_width_ftd_5 : STD_LOGIC;
  SIGNAL reg_out_width_ftd_6 : STD_LOGIC;
  SIGNAL nand_ssc : STD_LOGIC;
  SIGNAL reg_out_height_ftd : STD_LOGIC;
  SIGNAL reg_out_height_ftd_1 : STD_LOGIC;
  SIGNAL reg_out_height_ftd_2 : STD_LOGIC;
  SIGNAL reg_out_height_ftd_3 : STD_LOGIC;
  SIGNAL reg_out_height_ftd_4 : STD_LOGIC;
  SIGNAL reg_out_height_ftd_5 : STD_LOGIC;
  SIGNAL reg_out_height_ftd_6 : STD_LOGIC;

  SIGNAL and_58_nl : STD_LOGIC;
  SIGNAL max_val_and_nl : STD_LOGIC;
  SIGNAL not_73_nl : STD_LOGIC;
  SIGNAL LOOP_Y_mux_4_nl : STD_LOGIC;
  SIGNAL LOOP_Y_aelse_LOOP_Y_aelse_and_nl : STD_LOGIC;
  SIGNAL LOOP_WIDTH_acc_7_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LOOP_Y_acc_1_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL LOOP_Y_if_mul_5_nl : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL LOOP_Y_if_mux_5_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL LOOP_Y_else_acc_7_nl : STD_LOGIC_VECTOR (9 DOWNTO 0);
  SIGNAL and_146_nl : STD_LOGIC;
  SIGNAL LOOP_Y_if_mux_6_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL LOOP_CH_acc_2_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LOOP_CH_acc_3_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LOOP_HEIGHT_acc_2_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LOOP_HEIGHT_acc_3_nl : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL LOOP_X_acc_2_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL LOOP_X_acc_3_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL LOOP_Y_else_if_acc_nl : STD_LOGIC_VECTOR (12 DOWNTO 0);
  SIGNAL LOOP_Y_acc_2_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL LOOP_Y_if_LOOP_Y_if_and_1_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  SIGNAL LOOP_Y_if_mux_7_nl : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL LOOP_Y_if_mux_8_nl : STD_LOGIC_VECTOR (6 DOWNTO 0);
  COMPONENT UNET_IP_maxpool_run_max_run_max_fsm
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      arst_n : IN STD_LOGIC;
      fsm_output : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
      main_C_1_tr0 : IN STD_LOGIC;
      LOOP_CH_C_0_tr0 : IN STD_LOGIC;
      LOOP_HEIGHT_C_0_tr0 : IN STD_LOGIC;
      LOOP_WIDTH_C_0_tr0 : IN STD_LOGIC;
      LOOP_Y_C_0_tr0 : IN STD_LOGIC;
      LOOP_X_C_0_tr0 : IN STD_LOGIC;
      LOOP_WIDTH_C_3_tr0 : IN STD_LOGIC;
      LOOP_HEIGHT_C_1_tr0 : IN STD_LOGIC;
      LOOP_CH_C_1_tr0 : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL UNET_IP_maxpool_run_max_run_max_fsm_inst_fsm_output : STD_LOGIC_VECTOR (12
      DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0 : STD_LOGIC;
  SIGNAL UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0 : STD_LOGIC;

  FUNCTION CONV_SL_1_1(input_val:BOOLEAN)
  RETURN STD_LOGIC IS
  BEGIN
    IF input_val THEN RETURN '1';ELSE RETURN '0';END IF;
  END;

  FUNCTION MUX_s_1_2_2(input_0 : STD_LOGIC;
  input_1 : STD_LOGIC;
  sel : STD_LOGIC)
  RETURN STD_LOGIC IS
    VARIABLE result : STD_LOGIC;

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_10_2_2(input_0 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(9 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(9 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_12_2_2(input_0 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(11 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_3_2_2(input_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(2 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_4_2_2(input_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(3 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_6_2_2(input_0 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(5 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(5 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION MUX_v_7_2_2(input_0 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  input_1 : STD_LOGIC_VECTOR(6 DOWNTO 0);
  sel : STD_LOGIC)
  RETURN STD_LOGIC_VECTOR IS
    VARIABLE result : STD_LOGIC_VECTOR(6 DOWNTO 0);

    BEGIN
      CASE sel IS
        WHEN '0' =>
          result := input_0;
        WHEN others =>
          result := input_1;
      END CASE;
    RETURN result;
  END;

  FUNCTION minimum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1<arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION maximum(arg1,arg2:INTEGER) RETURN INTEGER IS
  BEGIN
    IF(arg1>arg2)THEN
      RETURN arg1;
    ELSE
      RETURN arg2;
    END IF;
  END;

  FUNCTION READSLICE_1_8(input_val:STD_LOGIC_VECTOR(7 DOWNTO 0);index:INTEGER)
  RETURN STD_LOGIC IS
    CONSTANT min_sat_index:INTEGER:= maximum( index, 0 );
    CONSTANT sat_index:INTEGER:= minimum( min_sat_index, 7);
  BEGIN
    RETURN input_val(sat_index);
  END;

BEGIN
  input_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_input_triosy_obj_ld_cse,
      lz => input_triosy_lz
    );
  output_triosy_obj : work.mgc_io_sync_pkg_v2.mgc_io_sync_v2
    GENERIC MAP(
      valid => 0
      )
    PORT MAP(
      ld => reg_input_triosy_obj_ld_cse,
      lz => output_triosy_lz
    );
  UNET_IP_maxpool_run_max_run_max_fsm_inst : UNET_IP_maxpool_run_max_run_max_fsm
    PORT MAP(
      clk => clk,
      rst => rst,
      arst_n => arst_n,
      fsm_output => UNET_IP_maxpool_run_max_run_max_fsm_inst_fsm_output,
      main_C_1_tr0 => exit_LOOP_CH_sva_mx0,
      LOOP_CH_C_0_tr0 => exit_LOOP_HEIGHT_sva_mx0,
      LOOP_HEIGHT_C_0_tr0 => UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0,
      LOOP_WIDTH_C_0_tr0 => exit_LOOP_X_sva_mx0,
      LOOP_Y_C_0_tr0 => UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0,
      LOOP_X_C_0_tr0 => exit_LOOP_X_sva_mx0,
      LOOP_WIDTH_C_3_tr0 => LOOP_Y_stage_0,
      LOOP_HEIGHT_C_1_tr0 => exit_LOOP_HEIGHT_sva_mx0,
      LOOP_CH_C_1_tr0 => exit_LOOP_CH_sva_mx0
    );
  fsm_output <= UNET_IP_maxpool_run_max_run_max_fsm_inst_fsm_output;
  UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_HEIGHT_C_0_tr0 <= NOT (READSLICE_1_8(STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'(
      '1' & (NOT reg_out_width_ftd) & (NOT reg_out_width_ftd_1) & (NOT reg_out_width_ftd_2)
      & (NOT reg_out_width_ftd_3) & (NOT reg_out_width_ftd_4) & (NOT reg_out_width_ftd_5)
      & (NOT reg_out_width_ftd_6)) + UNSIGNED'( "00000001"), 8)), 7));
  UNET_IP_maxpool_run_max_run_max_fsm_inst_LOOP_Y_C_0_tr0 <= NOT(LOOP_Y_stage_0_3
      OR LOOP_Y_stage_0_2 OR LOOP_Y_stage_0);

  nor_13_cse <= NOT(LOOP_Y_else_if_acc_itm_12_1 OR LOOP_Y_land_lpi_6_dfm_3);
  or_23_cse <= (fsm_output(1)) OR (fsm_output(11));
  nand_ssc <= NOT(and_dcpl_20 AND (NOT (fsm_output(1))));
  x_or_cse <= (fsm_output(4)) OR (fsm_output(6));
  LOOP_CH_acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT channels))
      + UNSIGNED'( "00000001"), 8));
  LOOP_CH_acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & c_sva_2) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      channels), 7), 8) + UNSIGNED'( "00000001"), 8));
  exit_LOOP_CH_sva_mx0 <= MUX_s_1_2_2((NOT (LOOP_CH_acc_2_nl(7))), (NOT (LOOP_CH_acc_3_nl(7))),
      fsm_output(11));
  c_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(c_sva) + UNSIGNED'( "0000001"),
      7));
  LOOP_HEIGHT_acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( '1' & (NOT reg_out_height_ftd)
      & (NOT reg_out_height_ftd_1) & (NOT reg_out_height_ftd_2) & (NOT reg_out_height_ftd_3)
      & (NOT reg_out_height_ftd_4) & (NOT reg_out_height_ftd_5) & (NOT reg_out_height_ftd_6))
      + UNSIGNED'( "00000001"), 8));
  LOOP_HEIGHT_acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & i_sva_2)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( (NOT reg_out_height_ftd) & (NOT reg_out_height_ftd_1)
      & (NOT reg_out_height_ftd_2) & (NOT reg_out_height_ftd_3) & (NOT reg_out_height_ftd_4)
      & (NOT reg_out_height_ftd_5) & (NOT reg_out_height_ftd_6)), 7), 8) + UNSIGNED'(
      "00000001"), 8));
  exit_LOOP_HEIGHT_sva_mx0 <= MUX_s_1_2_2((NOT (LOOP_HEIGHT_acc_2_nl(7))), (NOT (LOOP_HEIGHT_acc_3_nl(7))),
      fsm_output(10));
  i_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(i_sva) + UNSIGNED'( "0000001"),
      7));
  j_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(j_sva) + UNSIGNED'( "0000001"),
      7));
  LOOP_X_acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & (NOT pool_size))
      + UNSIGNED'( "0001"), 4));
  LOOP_X_acc_3_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & x_sva_2) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      pool_size), 3), 4) + UNSIGNED'( "0001"), 4));
  exit_LOOP_X_sva_mx0 <= MUX_s_1_2_2((NOT (LOOP_X_acc_2_nl(3))), (NOT (LOOP_X_acc_3_nl(3))),
      fsm_output(6));
  x_sva_2 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(x_sva) + UNSIGNED'( "001"),
      3));
  LOOP_Y_if_mul_4_ncse_sva_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(j_sva)
      * UNSIGNED(stride)), 10));
  LOOP_Y_else_if_acc_nl <= STD_LOGIC_VECTOR(CONV_SIGNED(CONV_SIGNED(CONV_SIGNED(SIGNED(max_val_13_2_lpi_3),
      12), 13) - CONV_SIGNED(CONV_SIGNED(SIGNED(input_rsci_q_d), 12), 13), 13));
  LOOP_Y_else_if_acc_itm_12_1 <= LOOP_Y_else_if_acc_nl(12);
  and_dcpl_20 <= NOT((fsm_output(0)) OR (fsm_output(12)));
  or_dcpl_21 <= (fsm_output(9)) OR (fsm_output(6)) OR (fsm_output(8));
  LOOP_Y_acc_2_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & y_sva) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(NOT
      pool_size), 3), 4) + UNSIGNED'( "0001"), 4));
  LOOP_Y_acc_2_itm_3_1 <= LOOP_Y_acc_2_nl(3);
  input_rsci_radr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(reg_LOOP_Y_if_acc_4_itm_1_cse)
      + UNSIGNED(z_out_5), 15));
  input_rsci_re_d_pff <= (NOT exit_LOOP_Y_sva_st_2) AND LOOP_Y_stage_0_3 AND (fsm_output(5));
  output_rsci_d_d <= max_val_13_2_lpi_5;
  output_rsci_wadr_d <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(LOOP_WIDTH_acc_6_itm),
      14), 15) + UNSIGNED(z_out_5), 15));
  output_rsci_we_d_pff <= fsm_output(8);
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd <= z_out_6;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_1 <= z_out_5_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_2 <= z_out_4_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_3 <= z_out_3;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_4 <= z_out_2;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_5 <= z_out_1;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( and_dcpl_20 = '0' ) THEN
        reg_out_width_ftd_6 <= z_out_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((NOT((CONV_SL_1_1(fsm_output(9 DOWNTO 5)=STD_LOGIC_VECTOR'("00000")))
          OR ((nor_13_cse OR LOOP_Y_asn_3_itm_3 OR (NOT LOOP_Y_stage_0_4)) AND (fsm_output(5)))))
          OR (fsm_output(4))) = '1' ) THEN
        max_val_13_2_lpi_3 <= MUX_v_12_2_2(max_val_13_2_lpi_5, input_rsci_q_d, and_58_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk, arst_n)
  BEGIN
    IF ( arst_n = '0' ) THEN
      reg_input_triosy_obj_ld_cse <= '0';
      LOOP_Y_asn_3_itm_3 <= '0';
      LOOP_Y_land_lpi_6_dfm_3 <= '0';
      exit_LOOP_Y_sva_st_2 <= '0';
      exit_LOOP_Y_sva_st_1 <= '0';
      y_sva <= STD_LOGIC_VECTOR'( "000");
      LOOP_Y_stage_0_2 <= '0';
      LOOP_Y_stage_0_3 <= '0';
      LOOP_Y_stage_0_4 <= '0';
      LOOP_Y_land_lpi_6_dfm_2 <= '0';
      LOOP_Y_land_lpi_6_dfm_1 <= '0';
    ELSIF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        reg_input_triosy_obj_ld_cse <= '0';
        LOOP_Y_asn_3_itm_3 <= '0';
        LOOP_Y_land_lpi_6_dfm_3 <= '0';
        exit_LOOP_Y_sva_st_2 <= '0';
        exit_LOOP_Y_sva_st_1 <= '0';
        y_sva <= STD_LOGIC_VECTOR'( "000");
        LOOP_Y_stage_0_2 <= '0';
        LOOP_Y_stage_0_3 <= '0';
        LOOP_Y_stage_0_4 <= '0';
        LOOP_Y_land_lpi_6_dfm_2 <= '0';
        LOOP_Y_land_lpi_6_dfm_1 <= '0';
      ELSE
        reg_input_triosy_obj_ld_cse <= exit_LOOP_CH_sva_mx0 AND or_23_cse;
        LOOP_Y_asn_3_itm_3 <= exit_LOOP_Y_sva_st_2;
        LOOP_Y_land_lpi_6_dfm_3 <= LOOP_Y_land_lpi_6_dfm_2;
        exit_LOOP_Y_sva_st_2 <= exit_LOOP_Y_sva_st_1;
        exit_LOOP_Y_sva_st_1 <= NOT LOOP_Y_acc_2_itm_3_1;
        y_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(LOOP_Y_acc_1_nl),
            3)), (fsm_output(5)));
        LOOP_Y_stage_0_2 <= LOOP_Y_stage_0 AND (fsm_output(5));
        LOOP_Y_stage_0_3 <= LOOP_Y_stage_0_2 AND (fsm_output(5));
        LOOP_Y_stage_0_4 <= LOOP_Y_stage_0_3 AND (fsm_output(5));
        LOOP_Y_land_lpi_6_dfm_2 <= LOOP_Y_land_lpi_6_dfm_1;
        LOOP_Y_land_lpi_6_dfm_1 <= NOT(CONV_SL_1_1(y_sva/=STD_LOGIC_VECTOR'("000"))
            OR CONV_SL_1_1(x_sva/=STD_LOGIC_VECTOR'("000")));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( or_23_cse = '1' ) THEN
        c_sva <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), c_sva_2, (fsm_output(11)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( nand_ssc = '1' ) THEN
        reg_out_height_ftd <= z_out_6;
        reg_out_height_ftd_1 <= z_out_5_1;
        reg_out_height_ftd_2 <= z_out_4_1;
        reg_out_height_ftd_3 <= z_out_3;
        reg_out_height_ftd_4 <= z_out_2;
        reg_out_height_ftd_5 <= z_out_1;
        reg_out_height_ftd_6 <= z_out_0;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( ((fsm_output(10)) OR (fsm_output(2))) = '1' ) THEN
        i_sva <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), i_sva_2, (fsm_output(10)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_dcpl_21 OR (fsm_output(4)) OR (fsm_output(7)))) = '1' ) THEN
        max_val_13_2_lpi_5 <= MUX_v_12_2_2(max_val_13_2_lpi_3, input_rsci_q_d, max_val_and_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      IF ( (NOT(or_dcpl_21 OR CONV_SL_1_1(fsm_output(5 DOWNTO 4)/=STD_LOGIC_VECTOR'("00"))))
          = '1' ) THEN
        j_sva <= MUX_v_7_2_2(STD_LOGIC_VECTOR'("0000000"), j_sva_2, not_73_nl);
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk, arst_n)
  BEGIN
    IF ( arst_n = '0' ) THEN
      x_sva <= STD_LOGIC_VECTOR'( "000");
    ELSIF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        x_sva <= STD_LOGIC_VECTOR'( "000");
      ELSIF ( x_or_cse = '1' ) THEN
        x_sva <= MUX_v_3_2_2(STD_LOGIC_VECTOR'("000"), x_sva_2, (fsm_output(6)));
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk, arst_n)
  BEGIN
    IF ( arst_n = '0' ) THEN
      LOOP_Y_stage_0 <= '0';
    ELSIF clk'EVENT AND ( clk = '1' ) THEN
      IF (rst = '1') THEN
        LOOP_Y_stage_0 <= '0';
      ELSIF ( (x_or_cse OR (fsm_output(5)) OR (fsm_output(7))) = '1' ) THEN
        LOOP_Y_stage_0 <= LOOP_Y_mux_4_nl OR x_or_cse;
      END IF;
    END IF;
  END PROCESS;
  PROCESS (clk)
  BEGIN
    IF clk'EVENT AND ( clk = '1' ) THEN
      reg_LOOP_Y_if_acc_4_itm_1_cse <= STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(LOOP_Y_if_mul_5_nl),
          15) + CONV_UNSIGNED(UNSIGNED(LOOP_Y_if_mux_5_nl), 15), 15));
      LOOP_Y_else_asn_itm_1 <= y_sva;
      LOOP_Y_if_acc_2_itm_1 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_4(9
          DOWNTO 0)) + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(x_sva), 3), 10), 10));
      LOOP_WIDTH_mul_1_itm <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(c_sva)
          * UNSIGNED(LOOP_Y_if_mux_6_nl)), 14));
      LOOP_WIDTH_acc_6_itm <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(z_out_4) +
          CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(j_sva), 7), 14), 14));
    END IF;
  END PROCESS;
  and_58_nl <= (LOOP_Y_else_if_acc_itm_12_1 OR LOOP_Y_land_lpi_6_dfm_3) AND (NOT
      LOOP_Y_asn_3_itm_3) AND LOOP_Y_stage_0_4 AND (fsm_output(5));
  LOOP_Y_acc_1_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(y_sva) + UNSIGNED'(
      "001"), 3));
  max_val_and_nl <= (NOT((nor_13_cse OR LOOP_Y_asn_3_itm_3) AND LOOP_Y_stage_0_4))
      AND (fsm_output(5));
  not_73_nl <= NOT (fsm_output(3));
  LOOP_Y_aelse_LOOP_Y_aelse_and_nl <= LOOP_Y_stage_0 AND LOOP_Y_acc_2_itm_3_1;
  LOOP_WIDTH_acc_7_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED('1' & j_sva_2) +
      CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'( (NOT reg_out_width_ftd) & (NOT reg_out_width_ftd_1)
      & (NOT reg_out_width_ftd_2) & (NOT reg_out_width_ftd_3) & (NOT reg_out_width_ftd_4)
      & (NOT reg_out_width_ftd_5) & (NOT reg_out_width_ftd_6)), 7), 8) + UNSIGNED'(
      "00000001"), 8));
  LOOP_Y_mux_4_nl <= MUX_s_1_2_2(LOOP_Y_aelse_LOOP_Y_aelse_and_nl, (NOT (LOOP_WIDTH_acc_7_nl(7))),
      fsm_output(7));
  LOOP_Y_if_mul_5_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(LOOP_Y_if_acc_2_itm_1)
      * UNSIGNED(width)), 15));
  LOOP_Y_else_acc_7_nl <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(LOOP_Y_if_mul_4_ncse_sva_1)
      + CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED(LOOP_Y_else_asn_itm_1), 3), 10), 10));
  and_146_nl <= (NOT LOOP_Y_land_lpi_6_dfm_1) AND (fsm_output(5));
  LOOP_Y_if_mux_5_nl <= MUX_v_10_2_2(LOOP_Y_if_mul_4_ncse_sva_1, STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED(LOOP_Y_else_acc_7_nl),
      10)), and_146_nl);
  LOOP_Y_if_mux_6_nl <= MUX_v_7_2_2(height, STD_LOGIC_VECTOR'( reg_out_height_ftd
      & reg_out_height_ftd_1 & reg_out_height_ftd_2 & reg_out_height_ftd_3 & reg_out_height_ftd_4
      & reg_out_height_ftd_5 & reg_out_height_ftd_6), fsm_output(7));
  mgc_div_7_3_0_b0_line_26 : PROCESS (width, height, fsm_output, stride)
    -- Interconnect Declarations
    VARIABLE divmod6448_2_diff_1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_diff_2 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_diff_3 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_diff_4 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_diff_5 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_diff_6 : STD_LOGIC_VECTOR (3 DOWNTO 0);
    VARIABLE divmod6448_2_lbuf_8_3 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_8_4 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_8_5 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_8_6 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_7_2 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_7_3 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_7_4 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_7_5 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_7_6 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6_1 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6_2 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6_3 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6_4 : STD_LOGIC;
    VARIABLE slc_fsm_output_1_5_ssc : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_6_5 : STD_LOGIC;
    VARIABLE divmod6448_2_lbuf_5_0 : STD_LOGIC_VECTOR (5 DOWNTO 0);

    VARIABLE divmod6448_2_loop951_7_acc_1_nl : STD_LOGIC_VECTOR (3 DOWNTO 0);
  BEGIN
    slc_fsm_output_1_5_ssc := fsm_output(1);
    divmod6448_2_lbuf_5_0 := MUX_v_6_2_2((width(5 DOWNTO 0)), (height(5 DOWNTO 0)),
        slc_fsm_output_1_5_ssc);
    divmod6448_2_lbuf_6_5 := MUX_s_1_2_2((width(6)), (height(6)), slc_fsm_output_1_5_ssc);
    divmod6448_2_diff_1 := STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(divmod6448_2_lbuf_6_5,
        1), 1), 4) + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_1(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_6_5 := divmod6448_2_diff_1(0);
    END IF;
    divmod6448_2_lbuf_7_2 := divmod6448_2_lbuf_6_5;
    divmod6448_2_lbuf_6 := divmod6448_2_lbuf_5_0(5);
    divmod6448_2_diff_2 := STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
        divmod6448_2_lbuf_6_5 & (divmod6448_2_lbuf_5_0(5))), 2), 4) + UNSIGNED('1'
        & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_2(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_7_2 := divmod6448_2_diff_2(1);
      divmod6448_2_lbuf_6 := divmod6448_2_diff_2(0);
    END IF;
    divmod6448_2_lbuf_8_3 := divmod6448_2_lbuf_7_2;
    divmod6448_2_lbuf_7_3 := divmod6448_2_lbuf_6;
    divmod6448_2_lbuf_6_1 := divmod6448_2_lbuf_5_0(4);
    divmod6448_2_diff_3 := STD_LOGIC_VECTOR(CONV_UNSIGNED(CONV_UNSIGNED(CONV_UNSIGNED(UNSIGNED'(
        divmod6448_2_lbuf_7_2 & divmod6448_2_lbuf_6 & (divmod6448_2_lbuf_5_0(4))),
        3), 4) + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_3(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_7_3 := divmod6448_2_diff_3(1);
      divmod6448_2_lbuf_8_3 := divmod6448_2_diff_3(2);
      divmod6448_2_lbuf_6_1 := divmod6448_2_diff_3(0);
    END IF;
    divmod6448_2_lbuf_8_4 := divmod6448_2_lbuf_7_3;
    divmod6448_2_lbuf_7_4 := divmod6448_2_lbuf_6_1;
    divmod6448_2_lbuf_6_2 := divmod6448_2_lbuf_5_0(3);
    divmod6448_2_diff_4 := STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( divmod6448_2_lbuf_8_3
        & divmod6448_2_lbuf_7_3 & divmod6448_2_lbuf_6_1 & (divmod6448_2_lbuf_5_0(3)))
        + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_4(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_7_4 := divmod6448_2_diff_4(1);
      divmod6448_2_lbuf_8_4 := divmod6448_2_diff_4(2);
      divmod6448_2_lbuf_6_2 := divmod6448_2_diff_4(0);
    END IF;
    divmod6448_2_lbuf_8_5 := divmod6448_2_lbuf_7_4;
    divmod6448_2_lbuf_7_5 := divmod6448_2_lbuf_6_2;
    divmod6448_2_lbuf_6_3 := divmod6448_2_lbuf_5_0(2);
    divmod6448_2_diff_5 := STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( divmod6448_2_lbuf_8_4
        & divmod6448_2_lbuf_7_4 & divmod6448_2_lbuf_6_2 & (divmod6448_2_lbuf_5_0(2)))
        + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_5(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_7_5 := divmod6448_2_diff_5(1);
      divmod6448_2_lbuf_8_5 := divmod6448_2_diff_5(2);
      divmod6448_2_lbuf_6_3 := divmod6448_2_diff_5(0);
    END IF;
    divmod6448_2_lbuf_8_6 := divmod6448_2_lbuf_7_5;
    divmod6448_2_lbuf_7_6 := divmod6448_2_lbuf_6_3;
    divmod6448_2_lbuf_6_4 := divmod6448_2_lbuf_5_0(1);
    divmod6448_2_diff_6 := STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( divmod6448_2_lbuf_8_5
        & divmod6448_2_lbuf_7_5 & divmod6448_2_lbuf_6_3 & (divmod6448_2_lbuf_5_0(1)))
        + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    IF ( (divmod6448_2_diff_6(3)) = '1' ) THEN
    ELSE
      divmod6448_2_lbuf_7_6 := divmod6448_2_diff_6(1);
      divmod6448_2_lbuf_8_6 := divmod6448_2_diff_6(2);
      divmod6448_2_lbuf_6_4 := divmod6448_2_diff_6(0);
    END IF;
    z_out_3 <= NOT (divmod6448_2_diff_4(3));
    z_out_2 <= NOT (divmod6448_2_diff_5(3));
    z_out_4_1 <= NOT (divmod6448_2_diff_3(3));
    z_out_1 <= NOT (divmod6448_2_diff_6(3));
    z_out_5_1 <= NOT (divmod6448_2_diff_2(3));
    divmod6448_2_loop951_7_acc_1_nl := STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'(
        divmod6448_2_lbuf_8_6 & divmod6448_2_lbuf_7_6 & divmod6448_2_lbuf_6_4 & (divmod6448_2_lbuf_5_0(0)))
        + UNSIGNED('1' & (NOT stride)) + UNSIGNED'( "0001"), 4));
    z_out_0 <= NOT (divmod6448_2_loop951_7_acc_1_nl(3));
    z_out_6 <= NOT (divmod6448_2_diff_1(3));
  END PROCESS mgc_div_7_3_0_b0_line_26;

  LOOP_Y_if_LOOP_Y_if_and_1_nl <= MUX_v_4_2_2(STD_LOGIC_VECTOR'("0000"), STD_LOGIC_VECTOR'(
      reg_out_width_ftd & reg_out_width_ftd_1 & reg_out_width_ftd_2 & reg_out_width_ftd_3),
      (fsm_output(7)));
  LOOP_Y_if_mux_7_nl <= MUX_v_3_2_2(stride, STD_LOGIC_VECTOR'( reg_out_width_ftd_4
      & reg_out_width_ftd_5 & reg_out_width_ftd_6), fsm_output(7));
  z_out_4 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(i_sva) * UNSIGNED(LOOP_Y_if_LOOP_Y_if_and_1_nl
      & LOOP_Y_if_mux_7_nl)), 14));
  LOOP_Y_if_mux_8_nl <= MUX_v_7_2_2(width, STD_LOGIC_VECTOR'( reg_out_width_ftd &
      reg_out_width_ftd_1 & reg_out_width_ftd_2 & reg_out_width_ftd_3 & reg_out_width_ftd_4
      & reg_out_width_ftd_5 & reg_out_width_ftd_6), fsm_output(8));
  z_out_5 <= STD_LOGIC_VECTOR(CONV_UNSIGNED(UNSIGNED'( UNSIGNED(LOOP_Y_if_mux_8_nl)
      * UNSIGNED(LOOP_WIDTH_mul_1_itm)), 15));
END v1;

-- ------------------------------------------------------------------
--  Design Unit:    UNET_IP_maxpool
-- ------------------------------------------------------------------

LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

USE work.mgc_io_sync_pkg_v2.ALL;


ENTITY UNET_IP_maxpool IS
  PORT(
    clk : IN STD_LOGIC;
    rst : IN STD_LOGIC;
    arst_n : IN STD_LOGIC;
    input_rsc_radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    input_rsc_re : OUT STD_LOGIC;
    input_rsc_q : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
    input_rsc_clken : OUT STD_LOGIC;
    input_triosy_lz : OUT STD_LOGIC;
    output_rsc_wadr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
    output_rsc_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
    output_rsc_we : OUT STD_LOGIC;
    output_rsc_clken : OUT STD_LOGIC;
    output_triosy_lz : OUT STD_LOGIC;
    channels : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    height : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    width : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
    pool_size : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
    stride : IN STD_LOGIC_VECTOR (2 DOWNTO 0)
  );
END UNET_IP_maxpool;

ARCHITECTURE v1 OF UNET_IP_maxpool IS
  -- Default Constants
  CONSTANT PWR : STD_LOGIC := '1';

  -- Interconnect Declarations
  SIGNAL input_rsci_q_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL input_rsci_radr_d : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL output_rsci_d_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL output_rsci_wadr_d : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL input_rsci_re_d_iff : STD_LOGIC;
  SIGNAL output_rsci_we_d_iff : STD_LOGIC;

  COMPONENT UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      q : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      re : OUT STD_LOGIC;
      radr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      q_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      radr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
      re_d : IN STD_LOGIC;
      readA_r_ram_ir_internal_RMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL input_rsci_q : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL input_rsci_radr : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL input_rsci_q_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL input_rsci_radr_d_1 : STD_LOGIC_VECTOR (14 DOWNTO 0);

  COMPONENT UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
    PORT(
      clken : OUT STD_LOGIC;
      we : OUT STD_LOGIC;
      d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      wadr : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      clken_d : IN STD_LOGIC;
      d_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      wadr_d : IN STD_LOGIC_VECTOR (14 DOWNTO 0);
      we_d : IN STD_LOGIC;
      writeA_w_ram_ir_internal_WMASK_B_d : IN STD_LOGIC
    );
  END COMPONENT;
  SIGNAL output_rsci_d : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL output_rsci_wadr : STD_LOGIC_VECTOR (14 DOWNTO 0);
  SIGNAL output_rsci_d_d_1 : STD_LOGIC_VECTOR (11 DOWNTO 0);
  SIGNAL output_rsci_wadr_d_1 : STD_LOGIC_VECTOR (14 DOWNTO 0);

  COMPONENT UNET_IP_maxpool_run_max
    PORT(
      clk : IN STD_LOGIC;
      rst : IN STD_LOGIC;
      arst_n : IN STD_LOGIC;
      input_triosy_lz : OUT STD_LOGIC;
      output_triosy_lz : OUT STD_LOGIC;
      channels : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
      height : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
      width : IN STD_LOGIC_VECTOR (6 DOWNTO 0);
      pool_size : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      stride : IN STD_LOGIC_VECTOR (2 DOWNTO 0);
      input_rsci_q_d : IN STD_LOGIC_VECTOR (11 DOWNTO 0);
      input_rsci_radr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      output_rsci_d_d : OUT STD_LOGIC_VECTOR (11 DOWNTO 0);
      output_rsci_wadr_d : OUT STD_LOGIC_VECTOR (14 DOWNTO 0);
      input_rsci_re_d_pff : OUT STD_LOGIC;
      output_rsci_we_d_pff : OUT STD_LOGIC
    );
  END COMPONENT;
  SIGNAL UNET_IP_maxpool_run_max_inst_channels : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_inst_height : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_inst_width : STD_LOGIC_VECTOR (6 DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_inst_pool_size : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_inst_stride : STD_LOGIC_VECTOR (2 DOWNTO 0);
  SIGNAL UNET_IP_maxpool_run_max_inst_input_rsci_q_d : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL UNET_IP_maxpool_run_max_inst_input_rsci_radr_d : STD_LOGIC_VECTOR (14 DOWNTO
      0);
  SIGNAL UNET_IP_maxpool_run_max_inst_output_rsci_d_d : STD_LOGIC_VECTOR (11 DOWNTO
      0);
  SIGNAL UNET_IP_maxpool_run_max_inst_output_rsci_wadr_d : STD_LOGIC_VECTOR (14 DOWNTO
      0);

BEGIN
  input_rsci : UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_rport_en_1_15_12_32768_1_32768_12_1_gen
    PORT MAP(
      clken => input_rsc_clken,
      q => input_rsci_q,
      re => input_rsc_re,
      radr => input_rsci_radr,
      clken_d => '1',
      q_d => input_rsci_q_d_1,
      radr_d => input_rsci_radr_d_1,
      re_d => input_rsci_re_d_iff,
      readA_r_ram_ir_internal_RMASK_B_d => input_rsci_re_d_iff
    );
  input_rsci_q <= input_rsc_q;
  input_rsc_radr <= input_rsci_radr;
  input_rsci_q_d <= input_rsci_q_d_1;
  input_rsci_radr_d_1 <= input_rsci_radr_d;

  output_rsci : UNET_IP_maxpool_Xilinx_RAMS_BLOCK_1R1W_RBW_wport_en_2_15_12_32768_1_32768_12_1_gen
    PORT MAP(
      clken => output_rsc_clken,
      we => output_rsc_we,
      d => output_rsci_d,
      wadr => output_rsci_wadr,
      clken_d => '1',
      d_d => output_rsci_d_d_1,
      wadr_d => output_rsci_wadr_d_1,
      we_d => output_rsci_we_d_iff,
      writeA_w_ram_ir_internal_WMASK_B_d => output_rsci_we_d_iff
    );
  output_rsc_d <= output_rsci_d;
  output_rsc_wadr <= output_rsci_wadr;
  output_rsci_d_d_1 <= output_rsci_d_d;
  output_rsci_wadr_d_1 <= output_rsci_wadr_d;

  UNET_IP_maxpool_run_max_inst : UNET_IP_maxpool_run_max
    PORT MAP(
      clk => clk,
      rst => rst,
      arst_n => arst_n,
      input_triosy_lz => input_triosy_lz,
      output_triosy_lz => output_triosy_lz,
      channels => UNET_IP_maxpool_run_max_inst_channels,
      height => UNET_IP_maxpool_run_max_inst_height,
      width => UNET_IP_maxpool_run_max_inst_width,
      pool_size => UNET_IP_maxpool_run_max_inst_pool_size,
      stride => UNET_IP_maxpool_run_max_inst_stride,
      input_rsci_q_d => UNET_IP_maxpool_run_max_inst_input_rsci_q_d,
      input_rsci_radr_d => UNET_IP_maxpool_run_max_inst_input_rsci_radr_d,
      output_rsci_d_d => UNET_IP_maxpool_run_max_inst_output_rsci_d_d,
      output_rsci_wadr_d => UNET_IP_maxpool_run_max_inst_output_rsci_wadr_d,
      input_rsci_re_d_pff => input_rsci_re_d_iff,
      output_rsci_we_d_pff => output_rsci_we_d_iff
    );
  UNET_IP_maxpool_run_max_inst_channels <= channels;
  UNET_IP_maxpool_run_max_inst_height <= height;
  UNET_IP_maxpool_run_max_inst_width <= width;
  UNET_IP_maxpool_run_max_inst_pool_size <= pool_size;
  UNET_IP_maxpool_run_max_inst_stride <= stride;
  UNET_IP_maxpool_run_max_inst_input_rsci_q_d <= input_rsci_q_d;
  input_rsci_radr_d <= UNET_IP_maxpool_run_max_inst_input_rsci_radr_d;
  output_rsci_d_d <= UNET_IP_maxpool_run_max_inst_output_rsci_d_d;
  output_rsci_wadr_d <= UNET_IP_maxpool_run_max_inst_output_rsci_wadr_d;

END v1;



